../hazard3/hdl/hazard3_config_inst.vh