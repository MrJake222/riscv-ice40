../hazard3_ops.vh