../hazard3/hdl/rv_opcodes.vh