../hazard3/hdl/hazard3_width_const.vh