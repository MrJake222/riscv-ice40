`define __ENABLE_FPU__
