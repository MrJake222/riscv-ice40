../configsoc.vh