../hazard3_config_inst.vh