../config.vh