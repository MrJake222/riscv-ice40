../rv_opcodes.vh