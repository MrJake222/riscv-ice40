../hazard3_csr_addr.vh