../hazard3/hdl/hazard3_csr_addr.vh