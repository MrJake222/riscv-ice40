`timescale 1 ns / 1 ns

module t20_custom ();

`include "dep.v"

initial
begin
	force soc.cpu_n_reset = 0;
	force soc.dbg_mem_op = 1'b1;
	force soc.dbg_wren = 4'hF;
	
    // Try to use stack
    // EXPECTED: stack ptr loaded with 10000 and decremented to FFF0
    //           x10 loads 20088 and saves it to stack address FFFC
    //           x11 is loaded from stack with 20088

    // program rom
force soc.dbg_adr = 32'h20000; force soc.dbg_do = 32'h00010137; #1000;
force soc.dbg_adr = 32'h20004; force soc.dbg_do = 32'h000036b7; #1000;
force soc.dbg_adr = 32'h20008; force soc.dbg_do = 32'h00000713; #1000;
force soc.dbg_adr = 32'h2000c; force soc.dbg_do = 32'hc0c68693; #1000;
force soc.dbg_adr = 32'h20010; force soc.dbg_do = 32'h02d77463; #1000;
force soc.dbg_adr = 32'h20014; force soc.dbg_do = 32'hfff68693; #1000;
force soc.dbg_adr = 32'h20018; force soc.dbg_do = 32'h40e686b3; #1000;
force soc.dbg_adr = 32'h2001c; force soc.dbg_do = 32'hffc6f693; #1000;
force soc.dbg_adr = 32'h20020; force soc.dbg_do = 32'h00468693; #1000;
force soc.dbg_adr = 32'h20024; force soc.dbg_do = 32'h00d70733; #1000;
force soc.dbg_adr = 32'h20028; force soc.dbg_do = 32'h00000793; #1000;
force soc.dbg_adr = 32'h2002c; force soc.dbg_do = 32'h00478793; #1000;
force soc.dbg_adr = 32'h20030; force soc.dbg_do = 32'hfe07ae23; #1000;
force soc.dbg_adr = 32'h20034; force soc.dbg_do = 32'hfee79ce3; #1000;
force soc.dbg_adr = 32'h20038; force soc.dbg_do = 32'h1240006f; #1000;
force soc.dbg_adr = 32'h2003c; force soc.dbg_do = 32'h00a00793; #1000;
force soc.dbg_adr = 32'h20040; force soc.dbg_do = 32'h02f50263; #1000;
force soc.dbg_adr = 32'h20044; force soc.dbg_do = 32'h00010737; #1000;
force soc.dbg_adr = 32'h20048; force soc.dbg_do = 32'h01470713; #1000;
force soc.dbg_adr = 32'h2004c; force soc.dbg_do = 32'h00072783; #1000;
force soc.dbg_adr = 32'h20050; force soc.dbg_do = 32'h0027f793; #1000;
force soc.dbg_adr = 32'h20054; force soc.dbg_do = 32'hfe078ce3; #1000;
force soc.dbg_adr = 32'h20058; force soc.dbg_do = 32'h000107b7; #1000;
force soc.dbg_adr = 32'h2005c; force soc.dbg_do = 32'h00a7a823; #1000;
force soc.dbg_adr = 32'h20060; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20064; force soc.dbg_do = 32'h00010737; #1000;
force soc.dbg_adr = 32'h20068; force soc.dbg_do = 32'h01470713; #1000;
force soc.dbg_adr = 32'h2006c; force soc.dbg_do = 32'h00072783; #1000;
force soc.dbg_adr = 32'h20070; force soc.dbg_do = 32'h0027f793; #1000;
force soc.dbg_adr = 32'h20074; force soc.dbg_do = 32'hfe078ce3; #1000;
force soc.dbg_adr = 32'h20078; force soc.dbg_do = 32'h000107b7; #1000;
force soc.dbg_adr = 32'h2007c; force soc.dbg_do = 32'h00d00713; #1000;
force soc.dbg_adr = 32'h20080; force soc.dbg_do = 32'h00e7a823; #1000;
force soc.dbg_adr = 32'h20084; force soc.dbg_do = 32'hfc1ff06f; #1000;
force soc.dbg_adr = 32'h20088; force soc.dbg_do = 32'hff010113; #1000;
force soc.dbg_adr = 32'h2008c; force soc.dbg_do = 32'h00058793; #1000;
force soc.dbg_adr = 32'h20090; force soc.dbg_do = 32'h00812423; #1000;
force soc.dbg_adr = 32'h20094; force soc.dbg_do = 32'h00a00593; #1000;
force soc.dbg_adr = 32'h20098; force soc.dbg_do = 32'h00050413; #1000;
force soc.dbg_adr = 32'h2009c; force soc.dbg_do = 32'h00078513; #1000;
force soc.dbg_adr = 32'h200a0; force soc.dbg_do = 32'h00112623; #1000;
force soc.dbg_adr = 32'h200a4; force soc.dbg_do = 32'h00912223; #1000;
force soc.dbg_adr = 32'h200a8; force soc.dbg_do = 32'h1cd030ef; #1000;
force soc.dbg_adr = 32'h200ac; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h200b0; force soc.dbg_do = 32'h00040513; #1000;
force soc.dbg_adr = 32'h200b4; force soc.dbg_do = 32'h1c1030ef; #1000;
force soc.dbg_adr = 32'h200b8; force soc.dbg_do = 32'h00a00593; #1000;
force soc.dbg_adr = 32'h200bc; force soc.dbg_do = 32'h00050493; #1000;
force soc.dbg_adr = 32'h200c0; force soc.dbg_do = 32'h1b5030ef; #1000;
force soc.dbg_adr = 32'h200c4; force soc.dbg_do = 32'h00050413; #1000;
force soc.dbg_adr = 32'h200c8; force soc.dbg_do = 32'h00a00593; #1000;
force soc.dbg_adr = 32'h200cc; force soc.dbg_do = 32'h00048513; #1000;
force soc.dbg_adr = 32'h200d0; force soc.dbg_do = 32'h229030ef; #1000;
force soc.dbg_adr = 32'h200d4; force soc.dbg_do = 32'h00400793; #1000;
force soc.dbg_adr = 32'h200d8; force soc.dbg_do = 32'h00a7a533; #1000;
force soc.dbg_adr = 32'h200dc; force soc.dbg_do = 32'h00c12083; #1000;
force soc.dbg_adr = 32'h200e0; force soc.dbg_do = 32'h00a40533; #1000;
force soc.dbg_adr = 32'h200e4; force soc.dbg_do = 32'h00812403; #1000;
force soc.dbg_adr = 32'h200e8; force soc.dbg_do = 32'h00412483; #1000;
force soc.dbg_adr = 32'h200ec; force soc.dbg_do = 32'h01010113; #1000;
force soc.dbg_adr = 32'h200f0; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h200f4; force soc.dbg_do = 32'hc0002573; #1000;
force soc.dbg_adr = 32'h200f8; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h200fc; force soc.dbg_do = 32'hc0202573; #1000;
force soc.dbg_adr = 32'h20100; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20104; force soc.dbg_do = 32'hc0002773; #1000;
force soc.dbg_adr = 32'h20108; force soc.dbg_do = 32'h000037b7; #1000;
force soc.dbg_adr = 32'h2010c; force soc.dbg_do = 32'hbee7a623; #1000;
force soc.dbg_adr = 32'h20110; force soc.dbg_do = 32'hc02026f3; #1000;
force soc.dbg_adr = 32'h20114; force soc.dbg_do = 32'h00003737; #1000;
force soc.dbg_adr = 32'h20118; force soc.dbg_do = 32'h000107b7; #1000;
force soc.dbg_adr = 32'h2011c; force soc.dbg_do = 32'hbed72423; #1000;
force soc.dbg_adr = 32'h20120; force soc.dbg_do = 32'h0187a703; #1000;
force soc.dbg_adr = 32'h20124; force soc.dbg_do = 32'h000037b7; #1000;
force soc.dbg_adr = 32'h20128; force soc.dbg_do = 32'hbee7a223; #1000;
force soc.dbg_adr = 32'h2012c; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20130; force soc.dbg_do = 32'hc0002773; #1000;
force soc.dbg_adr = 32'h20134; force soc.dbg_do = 32'h000037b7; #1000;
force soc.dbg_adr = 32'h20138; force soc.dbg_do = 32'hbee7a023; #1000;
force soc.dbg_adr = 32'h2013c; force soc.dbg_do = 32'hc02026f3; #1000;
force soc.dbg_adr = 32'h20140; force soc.dbg_do = 32'h00003737; #1000;
force soc.dbg_adr = 32'h20144; force soc.dbg_do = 32'h000107b7; #1000;
force soc.dbg_adr = 32'h20148; force soc.dbg_do = 32'hbcd72e23; #1000;
force soc.dbg_adr = 32'h2014c; force soc.dbg_do = 32'h0187a703; #1000;
force soc.dbg_adr = 32'h20150; force soc.dbg_do = 32'h000037b7; #1000;
force soc.dbg_adr = 32'h20154; force soc.dbg_do = 32'hbce7ac23; #1000;
force soc.dbg_adr = 32'h20158; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h2015c; force soc.dbg_do = 32'hfd010113; #1000;
force soc.dbg_adr = 32'h20160; force soc.dbg_do = 32'h02812423; #1000;
force soc.dbg_adr = 32'h20164; force soc.dbg_do = 32'h02912223; #1000;
force soc.dbg_adr = 32'h20168; force soc.dbg_do = 32'h000034b7; #1000;
force soc.dbg_adr = 32'h2016c; force soc.dbg_do = 32'h02112623; #1000;
force soc.dbg_adr = 32'h20170; force soc.dbg_do = 32'h03212023; #1000;
force soc.dbg_adr = 32'h20174; force soc.dbg_do = 32'h01312e23; #1000;
force soc.dbg_adr = 32'h20178; force soc.dbg_do = 32'h01412c23; #1000;
force soc.dbg_adr = 32'h2017c; force soc.dbg_do = 32'h01512a23; #1000;
force soc.dbg_adr = 32'h20180; force soc.dbg_do = 32'h01612823; #1000;
force soc.dbg_adr = 32'h20184; force soc.dbg_do = 32'h01712623; #1000;
force soc.dbg_adr = 32'h20188; force soc.dbg_do = 32'h01812423; #1000;
force soc.dbg_adr = 32'h2018c; force soc.dbg_do = 32'h00000793; #1000;
force soc.dbg_adr = 32'h20190; force soc.dbg_do = 32'hc0c48493; #1000;
force soc.dbg_adr = 32'h20194; force soc.dbg_do = 32'h0297f263; #1000;
force soc.dbg_adr = 32'h20198; force soc.dbg_do = 32'h00000413; #1000;
force soc.dbg_adr = 32'h2019c; force soc.dbg_do = 32'h00024937; #1000;
force soc.dbg_adr = 32'h201a0; force soc.dbg_do = 32'h00042603; #1000;
force soc.dbg_adr = 32'h201a4; force soc.dbg_do = 32'h00040593; #1000;
force soc.dbg_adr = 32'h201a8; force soc.dbg_do = 32'hb7490513; #1000;
force soc.dbg_adr = 32'h201ac; force soc.dbg_do = 32'h40040413; #1000;
force soc.dbg_adr = 32'h201b0; force soc.dbg_do = 32'h368020ef; #1000;
force soc.dbg_adr = 32'h201b4; force soc.dbg_do = 32'hfe9466e3; #1000;
force soc.dbg_adr = 32'h201b8; force soc.dbg_do = 32'h00012537; #1000;
force soc.dbg_adr = 32'h201bc; force soc.dbg_do = 32'hb3450513; #1000;
force soc.dbg_adr = 32'h201c0; force soc.dbg_do = 32'h490000ef; #1000;
force soc.dbg_adr = 32'h201c4; force soc.dbg_do = 32'h00003637; #1000;
force soc.dbg_adr = 32'h201c8; force soc.dbg_do = 32'h00003537; #1000;
force soc.dbg_adr = 32'h201cc; force soc.dbg_do = 32'h000035b7; #1000;
force soc.dbg_adr = 32'h201d0; force soc.dbg_do = 32'h000036b7; #1000;
force soc.dbg_adr = 32'h201d4; force soc.dbg_do = 32'h00003737; #1000;
force soc.dbg_adr = 32'h201d8; force soc.dbg_do = 32'h000037b7; #1000;
force soc.dbg_adr = 32'h201dc; force soc.dbg_do = 32'hbe872703; #1000;
force soc.dbg_adr = 32'h201e0; force soc.dbg_do = 32'hbe47a783; #1000;
force soc.dbg_adr = 32'h201e4; force soc.dbg_do = 32'hbec6a683; #1000;
force soc.dbg_adr = 32'h201e8; force soc.dbg_do = 32'hbd862903; #1000;
force soc.dbg_adr = 32'h201ec; force soc.dbg_do = 32'hbe052483; #1000;
force soc.dbg_adr = 32'h201f0; force soc.dbg_do = 32'hbdc5a403; #1000;
force soc.dbg_adr = 32'h201f4; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h201f8; force soc.dbg_do = 32'h000125b7; #1000;
force soc.dbg_adr = 32'h201fc; force soc.dbg_do = 32'hb3458593; #1000;
force soc.dbg_adr = 32'h20200; force soc.dbg_do = 32'hb8050513; #1000;
force soc.dbg_adr = 32'h20204; force soc.dbg_do = 32'h40e40433; #1000;
force soc.dbg_adr = 32'h20208; force soc.dbg_do = 32'h40d484b3; #1000;
force soc.dbg_adr = 32'h2020c; force soc.dbg_do = 32'h40f90933; #1000;
force soc.dbg_adr = 32'h20210; force soc.dbg_do = 32'h308020ef; #1000;
force soc.dbg_adr = 32'h20214; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20218; force soc.dbg_do = 32'h00048593; #1000;
force soc.dbg_adr = 32'h2021c; force soc.dbg_do = 32'hb8c50513; #1000;
force soc.dbg_adr = 32'h20220; force soc.dbg_do = 32'h2f8020ef; #1000;
force soc.dbg_adr = 32'h20224; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20228; force soc.dbg_do = 32'h00040593; #1000;
force soc.dbg_adr = 32'h2022c; force soc.dbg_do = 32'hb9850513; #1000;
force soc.dbg_adr = 32'h20230; force soc.dbg_do = 32'h2e8020ef; #1000;
force soc.dbg_adr = 32'h20234; force soc.dbg_do = 32'h000f45b7; #1000;
force soc.dbg_adr = 32'h20238; force soc.dbg_do = 32'h00090513; #1000;
force soc.dbg_adr = 32'h2023c; force soc.dbg_do = 32'h24058593; #1000;
force soc.dbg_adr = 32'h20240; force soc.dbg_do = 32'h0b9030ef; #1000;
force soc.dbg_adr = 32'h20244; force soc.dbg_do = 32'h000f45b7; #1000;
force soc.dbg_adr = 32'h20248; force soc.dbg_do = 32'h00050993; #1000;
force soc.dbg_adr = 32'h2024c; force soc.dbg_do = 32'h24058593; #1000;
force soc.dbg_adr = 32'h20250; force soc.dbg_do = 32'h00090513; #1000;
force soc.dbg_adr = 32'h20254; force soc.dbg_do = 32'h021030ef; #1000;
force soc.dbg_adr = 32'h20258; force soc.dbg_do = 32'h00050613; #1000;
force soc.dbg_adr = 32'h2025c; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20260; force soc.dbg_do = 32'h00098693; #1000;
force soc.dbg_adr = 32'h20264; force soc.dbg_do = 32'h00090593; #1000;
force soc.dbg_adr = 32'h20268; force soc.dbg_do = 32'hba450513; #1000;
force soc.dbg_adr = 32'h2026c; force soc.dbg_do = 32'h2ac020ef; #1000;
force soc.dbg_adr = 32'h20270; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20274; force soc.dbg_do = 32'hbc450513; #1000;
force soc.dbg_adr = 32'h20278; force soc.dbg_do = 32'h2a0020ef; #1000;
force soc.dbg_adr = 32'h2027c; force soc.dbg_do = 32'h41f4d993; #1000;
force soc.dbg_adr = 32'h20280; force soc.dbg_do = 32'h01b4d713; #1000;
force soc.dbg_adr = 32'h20284; force soc.dbg_do = 32'h00549693; #1000;
force soc.dbg_adr = 32'h20288; force soc.dbg_do = 32'h00599793; #1000;
force soc.dbg_adr = 32'h2028c; force soc.dbg_do = 32'h00f767b3; #1000;
force soc.dbg_adr = 32'h20290; force soc.dbg_do = 32'h40968733; #1000;
force soc.dbg_adr = 32'h20294; force soc.dbg_do = 32'h00e6b6b3; #1000;
force soc.dbg_adr = 32'h20298; force soc.dbg_do = 32'h413787b3; #1000;
force soc.dbg_adr = 32'h2029c; force soc.dbg_do = 32'h40d787b3; #1000;
force soc.dbg_adr = 32'h202a0; force soc.dbg_do = 32'h00279793; #1000;
force soc.dbg_adr = 32'h202a4; force soc.dbg_do = 32'h01e75693; #1000;
force soc.dbg_adr = 32'h202a8; force soc.dbg_do = 32'h00271713; #1000;
force soc.dbg_adr = 32'h202ac; force soc.dbg_do = 32'h00970533; #1000;
force soc.dbg_adr = 32'h202b0; force soc.dbg_do = 32'h00f6e7b3; #1000;
force soc.dbg_adr = 32'h202b4; force soc.dbg_do = 32'h00e53733; #1000;
force soc.dbg_adr = 32'h202b8; force soc.dbg_do = 32'h013787b3; #1000;
force soc.dbg_adr = 32'h202bc; force soc.dbg_do = 32'h00f707b3; #1000;
force soc.dbg_adr = 32'h202c0; force soc.dbg_do = 32'h41f45a13; #1000;
force soc.dbg_adr = 32'h202c4; force soc.dbg_do = 32'h00379793; #1000;
force soc.dbg_adr = 32'h202c8; force soc.dbg_do = 32'h01d55593; #1000;
force soc.dbg_adr = 32'h202cc; force soc.dbg_do = 32'h00f5e5b3; #1000;
force soc.dbg_adr = 32'h202d0; force soc.dbg_do = 32'h000a0693; #1000;
force soc.dbg_adr = 32'h202d4; force soc.dbg_do = 32'h00040613; #1000;
force soc.dbg_adr = 32'h202d8; force soc.dbg_do = 32'h00351513; #1000;
force soc.dbg_adr = 32'h202dc; force soc.dbg_do = 32'h3e8020ef; #1000;
force soc.dbg_adr = 32'h202e0; force soc.dbg_do = 32'h3e800613; #1000;
force soc.dbg_adr = 32'h202e4; force soc.dbg_do = 32'h00000693; #1000;
force soc.dbg_adr = 32'h202e8; force soc.dbg_do = 32'h00050c13; #1000;
force soc.dbg_adr = 32'h202ec; force soc.dbg_do = 32'h00058b93; #1000;
force soc.dbg_adr = 32'h202f0; force soc.dbg_do = 32'h19d020ef; #1000;
force soc.dbg_adr = 32'h202f4; force soc.dbg_do = 32'h00058a93; #1000;
force soc.dbg_adr = 32'h202f8; force soc.dbg_do = 32'h00050b13; #1000;
force soc.dbg_adr = 32'h202fc; force soc.dbg_do = 32'h3e800613; #1000;
force soc.dbg_adr = 32'h20300; force soc.dbg_do = 32'h00000693; #1000;
force soc.dbg_adr = 32'h20304; force soc.dbg_do = 32'h000c0513; #1000;
force soc.dbg_adr = 32'h20308; force soc.dbg_do = 32'h000b8593; #1000;
force soc.dbg_adr = 32'h2030c; force soc.dbg_do = 32'h3b8020ef; #1000;
force soc.dbg_adr = 32'h20310; force soc.dbg_do = 32'h00050613; #1000;
force soc.dbg_adr = 32'h20314; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20318; force soc.dbg_do = 32'h00058693; #1000;
force soc.dbg_adr = 32'h2031c; force soc.dbg_do = 32'h000a8793; #1000;
force soc.dbg_adr = 32'h20320; force soc.dbg_do = 32'h000b0713; #1000;
force soc.dbg_adr = 32'h20324; force soc.dbg_do = 32'hbc850513; #1000;
force soc.dbg_adr = 32'h20328; force soc.dbg_do = 32'h1f0020ef; #1000;
force soc.dbg_adr = 32'h2032c; force soc.dbg_do = 32'h01b45713; #1000;
force soc.dbg_adr = 32'h20330; force soc.dbg_do = 32'h00541693; #1000;
force soc.dbg_adr = 32'h20334; force soc.dbg_do = 32'h005a1793; #1000;
force soc.dbg_adr = 32'h20338; force soc.dbg_do = 32'h00f767b3; #1000;
force soc.dbg_adr = 32'h2033c; force soc.dbg_do = 32'h40868733; #1000;
force soc.dbg_adr = 32'h20340; force soc.dbg_do = 32'h00e6b6b3; #1000;
force soc.dbg_adr = 32'h20344; force soc.dbg_do = 32'h414787b3; #1000;
force soc.dbg_adr = 32'h20348; force soc.dbg_do = 32'h40d787b3; #1000;
force soc.dbg_adr = 32'h2034c; force soc.dbg_do = 32'h00279793; #1000;
force soc.dbg_adr = 32'h20350; force soc.dbg_do = 32'h01e75693; #1000;
force soc.dbg_adr = 32'h20354; force soc.dbg_do = 32'h00271713; #1000;
force soc.dbg_adr = 32'h20358; force soc.dbg_do = 32'h00870533; #1000;
force soc.dbg_adr = 32'h2035c; force soc.dbg_do = 32'h00f6e7b3; #1000;
force soc.dbg_adr = 32'h20360; force soc.dbg_do = 32'h00e53733; #1000;
force soc.dbg_adr = 32'h20364; force soc.dbg_do = 32'h014787b3; #1000;
force soc.dbg_adr = 32'h20368; force soc.dbg_do = 32'h00f707b3; #1000;
force soc.dbg_adr = 32'h2036c; force soc.dbg_do = 32'h00379793; #1000;
force soc.dbg_adr = 32'h20370; force soc.dbg_do = 32'h01d55593; #1000;
force soc.dbg_adr = 32'h20374; force soc.dbg_do = 32'h00f5e5b3; #1000;
force soc.dbg_adr = 32'h20378; force soc.dbg_do = 32'h00098693; #1000;
force soc.dbg_adr = 32'h2037c; force soc.dbg_do = 32'h00048613; #1000;
force soc.dbg_adr = 32'h20380; force soc.dbg_do = 32'h00351513; #1000;
force soc.dbg_adr = 32'h20384; force soc.dbg_do = 32'h340020ef; #1000;
force soc.dbg_adr = 32'h20388; force soc.dbg_do = 32'h3e800613; #1000;
force soc.dbg_adr = 32'h2038c; force soc.dbg_do = 32'h00000693; #1000;
force soc.dbg_adr = 32'h20390; force soc.dbg_do = 32'h00050a93; #1000;
force soc.dbg_adr = 32'h20394; force soc.dbg_do = 32'h00058a13; #1000;
force soc.dbg_adr = 32'h20398; force soc.dbg_do = 32'h0f5020ef; #1000;
force soc.dbg_adr = 32'h2039c; force soc.dbg_do = 32'h00050993; #1000;
force soc.dbg_adr = 32'h203a0; force soc.dbg_do = 32'h00058413; #1000;
force soc.dbg_adr = 32'h203a4; force soc.dbg_do = 32'h3e800613; #1000;
force soc.dbg_adr = 32'h203a8; force soc.dbg_do = 32'h00000693; #1000;
force soc.dbg_adr = 32'h203ac; force soc.dbg_do = 32'h000a8513; #1000;
force soc.dbg_adr = 32'h203b0; force soc.dbg_do = 32'h000a0593; #1000;
force soc.dbg_adr = 32'h203b4; force soc.dbg_do = 32'h310020ef; #1000;
force soc.dbg_adr = 32'h203b8; force soc.dbg_do = 32'h00050613; #1000;
force soc.dbg_adr = 32'h203bc; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h203c0; force soc.dbg_do = 32'h00098713; #1000;
force soc.dbg_adr = 32'h203c4; force soc.dbg_do = 32'h00040793; #1000;
force soc.dbg_adr = 32'h203c8; force soc.dbg_do = 32'h00058693; #1000;
force soc.dbg_adr = 32'h203cc; force soc.dbg_do = 32'hbdc50513; #1000;
force soc.dbg_adr = 32'h203d0; force soc.dbg_do = 32'h148020ef; #1000;
force soc.dbg_adr = 32'h203d4; force soc.dbg_do = 32'h00090513; #1000;
force soc.dbg_adr = 32'h203d8; force soc.dbg_do = 32'h5c4030ef; #1000;
force soc.dbg_adr = 32'h203dc; force soc.dbg_do = 32'h000247b7; #1000;
force soc.dbg_adr = 32'h203e0; force soc.dbg_do = 32'h00058693; #1000;
force soc.dbg_adr = 32'h203e4; force soc.dbg_do = 32'h00050613; #1000;
force soc.dbg_adr = 32'h203e8; force soc.dbg_do = 32'h30c7a583; #1000;
force soc.dbg_adr = 32'h203ec; force soc.dbg_do = 32'h3087a503; #1000;
force soc.dbg_adr = 32'h203f0; force soc.dbg_do = 32'h56d020ef; #1000;
force soc.dbg_adr = 32'h203f4; force soc.dbg_do = 32'h52c030ef; #1000;
force soc.dbg_adr = 32'h203f8; force soc.dbg_do = 32'h3e800593; #1000;
force soc.dbg_adr = 32'h203fc; force soc.dbg_do = 32'h00050413; #1000;
force soc.dbg_adr = 32'h20400; force soc.dbg_do = 32'h67c030ef; #1000;
force soc.dbg_adr = 32'h20404; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h20408; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h2040c; force soc.dbg_do = 32'hbf050513; #1000;
force soc.dbg_adr = 32'h20410; force soc.dbg_do = 32'h108020ef; #1000;
force soc.dbg_adr = 32'h20414; force soc.dbg_do = 32'h00040513; #1000;
force soc.dbg_adr = 32'h20418; force soc.dbg_do = 32'h6dd00593; #1000;
force soc.dbg_adr = 32'h2041c; force soc.dbg_do = 32'h660030ef; #1000;
force soc.dbg_adr = 32'h20420; force soc.dbg_do = 32'h3e800593; #1000;
force soc.dbg_adr = 32'h20424; force soc.dbg_do = 32'h00050993; #1000;
force soc.dbg_adr = 32'h20428; force soc.dbg_do = 32'h69c030ef; #1000;
force soc.dbg_adr = 32'h2042c; force soc.dbg_do = 32'h00050413; #1000;
force soc.dbg_adr = 32'h20430; force soc.dbg_do = 32'h3e800593; #1000;
force soc.dbg_adr = 32'h20434; force soc.dbg_do = 32'h00098513; #1000;
force soc.dbg_adr = 32'h20438; force soc.dbg_do = 32'h644030ef; #1000;
force soc.dbg_adr = 32'h2043c; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h20440; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20444; force soc.dbg_do = 32'h00040613; #1000;
force soc.dbg_adr = 32'h20448; force soc.dbg_do = 32'hc0c50513; #1000;
force soc.dbg_adr = 32'h2044c; force soc.dbg_do = 32'h0cc020ef; #1000;
force soc.dbg_adr = 32'h20450; force soc.dbg_do = 32'h00090513; #1000;
force soc.dbg_adr = 32'h20454; force soc.dbg_do = 32'h00a00593; #1000;
force soc.dbg_adr = 32'h20458; force soc.dbg_do = 32'h61c030ef; #1000;
force soc.dbg_adr = 32'h2045c; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h20460; force soc.dbg_do = 32'h00048513; #1000;
force soc.dbg_adr = 32'h20464; force soc.dbg_do = 32'h610030ef; #1000;
force soc.dbg_adr = 32'h20468; force soc.dbg_do = 32'h00a00593; #1000;
force soc.dbg_adr = 32'h2046c; force soc.dbg_do = 32'h00050493; #1000;
force soc.dbg_adr = 32'h20470; force soc.dbg_do = 32'h604030ef; #1000;
force soc.dbg_adr = 32'h20474; force soc.dbg_do = 32'h00050413; #1000;
force soc.dbg_adr = 32'h20478; force soc.dbg_do = 32'h00a00593; #1000;
force soc.dbg_adr = 32'h2047c; force soc.dbg_do = 32'h00048513; #1000;
force soc.dbg_adr = 32'h20480; force soc.dbg_do = 32'h678030ef; #1000;
force soc.dbg_adr = 32'h20484; force soc.dbg_do = 32'h00400793; #1000;
force soc.dbg_adr = 32'h20488; force soc.dbg_do = 32'h00a7a7b3; #1000;
force soc.dbg_adr = 32'h2048c; force soc.dbg_do = 32'h00f40433; #1000;
force soc.dbg_adr = 32'h20490; force soc.dbg_do = 32'h00040593; #1000;
force soc.dbg_adr = 32'h20494; force soc.dbg_do = 32'h00098513; #1000;
force soc.dbg_adr = 32'h20498; force soc.dbg_do = 32'h5e4030ef; #1000;
force soc.dbg_adr = 32'h2049c; force soc.dbg_do = 32'h3e800593; #1000;
force soc.dbg_adr = 32'h204a0; force soc.dbg_do = 32'h00050913; #1000;
force soc.dbg_adr = 32'h204a4; force soc.dbg_do = 32'h654030ef; #1000;
force soc.dbg_adr = 32'h204a8; force soc.dbg_do = 32'h00050493; #1000;
force soc.dbg_adr = 32'h204ac; force soc.dbg_do = 32'h3e800593; #1000;
force soc.dbg_adr = 32'h204b0; force soc.dbg_do = 32'h00090513; #1000;
force soc.dbg_adr = 32'h204b4; force soc.dbg_do = 32'h5c0030ef; #1000;
force soc.dbg_adr = 32'h204b8; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h204bc; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h204c0; force soc.dbg_do = 32'h00040693; #1000;
force soc.dbg_adr = 32'h204c4; force soc.dbg_do = 32'h00048613; #1000;
force soc.dbg_adr = 32'h204c8; force soc.dbg_do = 32'hc1c50513; #1000;
force soc.dbg_adr = 32'h204cc; force soc.dbg_do = 32'h04c020ef; #1000;
force soc.dbg_adr = 32'h204d0; force soc.dbg_do = 32'h0000006f; #1000;
force soc.dbg_adr = 32'h204d4; force soc.dbg_do = 32'h00003637; #1000;
force soc.dbg_adr = 32'h204d8; force soc.dbg_do = 32'hc0462703; #1000;
force soc.dbg_adr = 32'h204dc; force soc.dbg_do = 32'h00052783; #1000;
force soc.dbg_adr = 32'h204e0; force soc.dbg_do = 32'h00072583; #1000;
force soc.dbg_adr = 32'h204e4; force soc.dbg_do = 32'h02c72683; #1000;
force soc.dbg_adr = 32'h204e8; force soc.dbg_do = 32'h00472383; #1000;
force soc.dbg_adr = 32'h204ec; force soc.dbg_do = 32'h00872283; #1000;
force soc.dbg_adr = 32'h204f0; force soc.dbg_do = 32'h01072f83; #1000;
force soc.dbg_adr = 32'h204f4; force soc.dbg_do = 32'h01472f03; #1000;
force soc.dbg_adr = 32'h204f8; force soc.dbg_do = 32'h01872e83; #1000;
force soc.dbg_adr = 32'h204fc; force soc.dbg_do = 32'h01c72e03; #1000;
force soc.dbg_adr = 32'h20500; force soc.dbg_do = 32'h02072303; #1000;
force soc.dbg_adr = 32'h20504; force soc.dbg_do = 32'h02472883; #1000;
force soc.dbg_adr = 32'h20508; force soc.dbg_do = 32'h02872803; #1000;
force soc.dbg_adr = 32'h2050c; force soc.dbg_do = 32'h00b7a023; #1000;
force soc.dbg_adr = 32'h20510; force soc.dbg_do = 32'h00052583; #1000;
force soc.dbg_adr = 32'h20514; force soc.dbg_do = 32'h02d7a623; #1000;
force soc.dbg_adr = 32'h20518; force soc.dbg_do = 32'h0077a223; #1000;
force soc.dbg_adr = 32'h2051c; force soc.dbg_do = 32'h00500693; #1000;
force soc.dbg_adr = 32'h20520; force soc.dbg_do = 32'h0057a423; #1000;
force soc.dbg_adr = 32'h20524; force soc.dbg_do = 32'h01f7a823; #1000;
force soc.dbg_adr = 32'h20528; force soc.dbg_do = 32'h01e7aa23; #1000;
force soc.dbg_adr = 32'h2052c; force soc.dbg_do = 32'h01d7ac23; #1000;
force soc.dbg_adr = 32'h20530; force soc.dbg_do = 32'h01c7ae23; #1000;
force soc.dbg_adr = 32'h20534; force soc.dbg_do = 32'h0267a023; #1000;
force soc.dbg_adr = 32'h20538; force soc.dbg_do = 32'h0317a223; #1000;
force soc.dbg_adr = 32'h2053c; force soc.dbg_do = 32'h0307a423; #1000;
force soc.dbg_adr = 32'h20540; force soc.dbg_do = 32'h00d52623; #1000;
force soc.dbg_adr = 32'h20544; force soc.dbg_do = 32'h00b7a023; #1000;
force soc.dbg_adr = 32'h20548; force soc.dbg_do = 32'h00072703; #1000;
force soc.dbg_adr = 32'h2054c; force soc.dbg_do = 32'h000035b7; #1000;
force soc.dbg_adr = 32'h20550; force soc.dbg_do = 32'hbfc5a583; #1000;
force soc.dbg_adr = 32'h20554; force soc.dbg_do = 32'h00e7a023; #1000;
force soc.dbg_adr = 32'h20558; force soc.dbg_do = 32'hc0462703; #1000;
force soc.dbg_adr = 32'h2055c; force soc.dbg_do = 32'h00d7a623; #1000;
force soc.dbg_adr = 32'h20560; force soc.dbg_do = 32'h00c58693; #1000;
force soc.dbg_adr = 32'h20564; force soc.dbg_do = 32'h00d72623; #1000;
force soc.dbg_adr = 32'h20568; force soc.dbg_do = 32'h0047a683; #1000;
force soc.dbg_adr = 32'h2056c; force soc.dbg_do = 32'h06068663; #1000;
force soc.dbg_adr = 32'h20570; force soc.dbg_do = 32'h00052783; #1000;
force soc.dbg_adr = 32'h20574; force soc.dbg_do = 32'h0007af83; #1000;
force soc.dbg_adr = 32'h20578; force soc.dbg_do = 32'h0047af03; #1000;
force soc.dbg_adr = 32'h2057c; force soc.dbg_do = 32'h0087ae83; #1000;
force soc.dbg_adr = 32'h20580; force soc.dbg_do = 32'h00c7ae03; #1000;
force soc.dbg_adr = 32'h20584; force soc.dbg_do = 32'h0107a303; #1000;
force soc.dbg_adr = 32'h20588; force soc.dbg_do = 32'h0147a883; #1000;
force soc.dbg_adr = 32'h2058c; force soc.dbg_do = 32'h0187a803; #1000;
force soc.dbg_adr = 32'h20590; force soc.dbg_do = 32'h01c7a583; #1000;
force soc.dbg_adr = 32'h20594; force soc.dbg_do = 32'h0207a603; #1000;
force soc.dbg_adr = 32'h20598; force soc.dbg_do = 32'h0247a683; #1000;
force soc.dbg_adr = 32'h2059c; force soc.dbg_do = 32'h0287a703; #1000;
force soc.dbg_adr = 32'h205a0; force soc.dbg_do = 32'h02c7a783; #1000;
force soc.dbg_adr = 32'h205a4; force soc.dbg_do = 32'h01f52023; #1000;
force soc.dbg_adr = 32'h205a8; force soc.dbg_do = 32'h01e52223; #1000;
force soc.dbg_adr = 32'h205ac; force soc.dbg_do = 32'h01d52423; #1000;
force soc.dbg_adr = 32'h205b0; force soc.dbg_do = 32'h01c52623; #1000;
force soc.dbg_adr = 32'h205b4; force soc.dbg_do = 32'h00652823; #1000;
force soc.dbg_adr = 32'h205b8; force soc.dbg_do = 32'h01152a23; #1000;
force soc.dbg_adr = 32'h205bc; force soc.dbg_do = 32'h01052c23; #1000;
force soc.dbg_adr = 32'h205c0; force soc.dbg_do = 32'h00b52e23; #1000;
force soc.dbg_adr = 32'h205c4; force soc.dbg_do = 32'h02c52023; #1000;
force soc.dbg_adr = 32'h205c8; force soc.dbg_do = 32'h02d52223; #1000;
force soc.dbg_adr = 32'h205cc; force soc.dbg_do = 32'h02e52423; #1000;
force soc.dbg_adr = 32'h205d0; force soc.dbg_do = 32'h02f52623; #1000;
force soc.dbg_adr = 32'h205d4; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h205d8; force soc.dbg_do = 32'h00852683; #1000;
force soc.dbg_adr = 32'h205dc; force soc.dbg_do = 32'h00600613; #1000;
force soc.dbg_adr = 32'h205e0; force soc.dbg_do = 32'h00c7a623; #1000;
force soc.dbg_adr = 32'h205e4; force soc.dbg_do = 32'h00200613; #1000;
force soc.dbg_adr = 32'h205e8; force soc.dbg_do = 32'h04c68263; #1000;
force soc.dbg_adr = 32'h205ec; force soc.dbg_do = 32'h00300513; #1000;
force soc.dbg_adr = 32'h205f0; force soc.dbg_do = 32'h00a7a423; #1000;
force soc.dbg_adr = 32'h205f4; force soc.dbg_do = 32'h00100513; #1000;
force soc.dbg_adr = 32'h205f8; force soc.dbg_do = 32'h02a68263; #1000;
force soc.dbg_adr = 32'h205fc; force soc.dbg_do = 32'h00400593; #1000;
force soc.dbg_adr = 32'h20600; force soc.dbg_do = 32'h04b68463; #1000;
force soc.dbg_adr = 32'h20604; force soc.dbg_do = 32'h02068063; #1000;
force soc.dbg_adr = 32'h20608; force soc.dbg_do = 32'h00072703; #1000;
force soc.dbg_adr = 32'h2060c; force soc.dbg_do = 32'h01200693; #1000;
force soc.dbg_adr = 32'h20610; force soc.dbg_do = 32'h00d7a623; #1000;
force soc.dbg_adr = 32'h20614; force soc.dbg_do = 32'h00e7a023; #1000;
force soc.dbg_adr = 32'h20618; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h2061c; force soc.dbg_do = 32'h06400693; #1000;
force soc.dbg_adr = 32'h20620; force soc.dbg_do = 32'hfeb6d4e3; #1000;
force soc.dbg_adr = 32'h20624; force soc.dbg_do = 32'h0007a423; #1000;
force soc.dbg_adr = 32'h20628; force soc.dbg_do = 32'hfe1ff06f; #1000;
force soc.dbg_adr = 32'h2062c; force soc.dbg_do = 32'h00072703; #1000;
force soc.dbg_adr = 32'h20630; force soc.dbg_do = 32'h00100693; #1000;
force soc.dbg_adr = 32'h20634; force soc.dbg_do = 32'h00d7a423; #1000;
force soc.dbg_adr = 32'h20638; force soc.dbg_do = 32'h01200693; #1000;
force soc.dbg_adr = 32'h2063c; force soc.dbg_do = 32'h00d7a623; #1000;
force soc.dbg_adr = 32'h20640; force soc.dbg_do = 32'h00e7a023; #1000;
force soc.dbg_adr = 32'h20644; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20648; force soc.dbg_do = 32'h00c7a423; #1000;
force soc.dbg_adr = 32'h2064c; force soc.dbg_do = 32'hfbdff06f; #1000;
force soc.dbg_adr = 32'h20650; force soc.dbg_do = 32'hf7010113; #1000;
force soc.dbg_adr = 32'h20654; force soc.dbg_do = 32'h00050713; #1000;
force soc.dbg_adr = 32'h20658; force soc.dbg_do = 32'h03000513; #1000;
force soc.dbg_adr = 32'h2065c; force soc.dbg_do = 32'h00d12423; #1000;
force soc.dbg_adr = 32'h20660; force soc.dbg_do = 32'h00f12023; #1000;
force soc.dbg_adr = 32'h20664; force soc.dbg_do = 32'h08112623; #1000;
force soc.dbg_adr = 32'h20668; force soc.dbg_do = 32'h08812423; #1000;
force soc.dbg_adr = 32'h2066c; force soc.dbg_do = 32'h07612823; #1000;
force soc.dbg_adr = 32'h20670; force soc.dbg_do = 32'h05b12e23; #1000;
force soc.dbg_adr = 32'h20674; force soc.dbg_do = 32'h00e12623; #1000;
force soc.dbg_adr = 32'h20678; force soc.dbg_do = 32'h08912223; #1000;
force soc.dbg_adr = 32'h2067c; force soc.dbg_do = 32'h09212023; #1000;
force soc.dbg_adr = 32'h20680; force soc.dbg_do = 32'h07312e23; #1000;
force soc.dbg_adr = 32'h20684; force soc.dbg_do = 32'h07412c23; #1000;
force soc.dbg_adr = 32'h20688; force soc.dbg_do = 32'h07512a23; #1000;
force soc.dbg_adr = 32'h2068c; force soc.dbg_do = 32'h07712623; #1000;
force soc.dbg_adr = 32'h20690; force soc.dbg_do = 32'h07812423; #1000;
force soc.dbg_adr = 32'h20694; force soc.dbg_do = 32'h07912223; #1000;
force soc.dbg_adr = 32'h20698; force soc.dbg_do = 32'h005000ef; #1000;
force soc.dbg_adr = 32'h2069c; force soc.dbg_do = 32'h00050713; #1000;
force soc.dbg_adr = 32'h206a0; force soc.dbg_do = 32'h00003437; #1000;
force soc.dbg_adr = 32'h206a4; force soc.dbg_do = 32'h03000513; #1000;
force soc.dbg_adr = 32'h206a8; force soc.dbg_do = 32'hc0e42023; #1000;
force soc.dbg_adr = 32'h206ac; force soc.dbg_do = 32'h7f0000ef; #1000;
force soc.dbg_adr = 32'h206b0; force soc.dbg_do = 32'hc0042803; #1000;
force soc.dbg_adr = 32'h206b4; force soc.dbg_do = 32'h00003b37; #1000;
force soc.dbg_adr = 32'h206b8; force soc.dbg_do = 32'h00200613; #1000;
force soc.dbg_adr = 32'h206bc; force soc.dbg_do = 32'h02800713; #1000;
force soc.dbg_adr = 32'h206c0; force soc.dbg_do = 32'hc0ab2223; #1000;
force soc.dbg_adr = 32'h206c4; force soc.dbg_do = 32'h000245b7; #1000;
force soc.dbg_adr = 32'h206c8; force soc.dbg_do = 32'h01052023; #1000;
force soc.dbg_adr = 32'h206cc; force soc.dbg_do = 32'h00c52423; #1000;
force soc.dbg_adr = 32'h206d0; force soc.dbg_do = 32'h00e52623; #1000;
force soc.dbg_adr = 32'h206d4; force soc.dbg_do = 32'h00052223; #1000;
force soc.dbg_adr = 32'h206d8; force soc.dbg_do = 32'hc3c58593; #1000;
force soc.dbg_adr = 32'h206dc; force soc.dbg_do = 32'h01050513; #1000;
force soc.dbg_adr = 32'h206e0; force soc.dbg_do = 32'h7e8000ef; #1000;
force soc.dbg_adr = 32'h206e4; force soc.dbg_do = 32'h000245b7; #1000;
force soc.dbg_adr = 32'h206e8; force soc.dbg_do = 32'hc5c58593; #1000;
force soc.dbg_adr = 32'h206ec; force soc.dbg_do = 32'h01010513; #1000;
force soc.dbg_adr = 32'h206f0; force soc.dbg_do = 32'h7d8000ef; #1000;
force soc.dbg_adr = 32'h206f4; force soc.dbg_do = 32'h00024437; #1000;
force soc.dbg_adr = 32'h206f8; force soc.dbg_do = 32'h00a00613; #1000;
force soc.dbg_adr = 32'h206fc; force soc.dbg_do = 32'h0c800d93; #1000;
force soc.dbg_adr = 32'h20700; force soc.dbg_do = 32'hbc440513; #1000;
force soc.dbg_adr = 32'h20704; force soc.dbg_do = 32'h64cdae23; #1000;
force soc.dbg_adr = 32'h20708; force soc.dbg_do = 32'h611010ef; #1000;
force soc.dbg_adr = 32'h2070c; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20710; force soc.dbg_do = 32'hc7c50513; #1000;
force soc.dbg_adr = 32'h20714; force soc.dbg_do = 32'h605010ef; #1000;
force soc.dbg_adr = 32'h20718; force soc.dbg_do = 32'hbc440513; #1000;
force soc.dbg_adr = 32'h2071c; force soc.dbg_do = 32'h5fd010ef; #1000;
force soc.dbg_adr = 32'h20720; force soc.dbg_do = 32'h00003637; #1000;
force soc.dbg_adr = 32'h20724; force soc.dbg_do = 32'hbf062603; #1000;
force soc.dbg_adr = 32'h20728; force soc.dbg_do = 32'h00012783; #1000;
force soc.dbg_adr = 32'h2072c; force soc.dbg_do = 32'h00812683; #1000;
force soc.dbg_adr = 32'h20730; force soc.dbg_do = 32'h52060863; #1000;
force soc.dbg_adr = 32'h20734; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20738; force soc.dbg_do = 32'hcac50513; #1000;
force soc.dbg_adr = 32'h2073c; force soc.dbg_do = 32'h5dd010ef; #1000;
force soc.dbg_adr = 32'h20740; force soc.dbg_do = 32'hbc440513; #1000;
force soc.dbg_adr = 32'h20744; force soc.dbg_do = 32'h5d5010ef; #1000;
force soc.dbg_adr = 32'h20748; force soc.dbg_do = 32'h00012783; #1000;
force soc.dbg_adr = 32'h2074c; force soc.dbg_do = 32'h00812683; #1000;
force soc.dbg_adr = 32'h20750; force soc.dbg_do = 32'h00c12403; #1000;
force soc.dbg_adr = 32'h20754; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20758; force soc.dbg_do = 32'hd0850513; #1000;
force soc.dbg_adr = 32'h2075c; force soc.dbg_do = 32'h00040593; #1000;
force soc.dbg_adr = 32'h20760; force soc.dbg_do = 32'h00d12423; #1000;
force soc.dbg_adr = 32'h20764; force soc.dbg_do = 32'h00f12023; #1000;
force soc.dbg_adr = 32'h20768; force soc.dbg_do = 32'h5b1010ef; #1000;
force soc.dbg_adr = 32'h2076c; force soc.dbg_do = 32'h999ff0ef; #1000;
force soc.dbg_adr = 32'h20770; force soc.dbg_do = 32'h00012783; #1000;
force soc.dbg_adr = 32'h20774; force soc.dbg_do = 32'h00812683; #1000;
force soc.dbg_adr = 32'h20778; force soc.dbg_do = 32'h50805a63; #1000;
force soc.dbg_adr = 32'h2077c; force soc.dbg_do = 32'h07a12023; #1000;
force soc.dbg_adr = 32'h20780; force soc.dbg_do = 32'h00100d13; #1000;
force soc.dbg_adr = 32'h20784; force soc.dbg_do = 32'h00001bb7; #1000;
force soc.dbg_adr = 32'h20788; force soc.dbg_do = 32'h000037b7; #1000;
force soc.dbg_adr = 32'h2078c; force soc.dbg_do = 32'h04300c93; #1000;
force soc.dbg_adr = 32'h20790; force soc.dbg_do = 32'h000d0c13; #1000;
force soc.dbg_adr = 32'h20794; force soc.dbg_do = 32'h00000413; #1000;
force soc.dbg_adr = 32'h20798; force soc.dbg_do = 32'h0c8b8b93; #1000;
force soc.dbg_adr = 32'h2079c; force soc.dbg_do = 32'h00f12023; #1000;
force soc.dbg_adr = 32'h207a0; force soc.dbg_do = 32'h00003ab7; #1000;
force soc.dbg_adr = 32'h207a4; force soc.dbg_do = 32'h000039b7; #1000;
force soc.dbg_adr = 32'h207a8; force soc.dbg_do = 32'h03010913; #1000;
force soc.dbg_adr = 32'h207ac; force soc.dbg_do = 32'h00003a37; #1000;
force soc.dbg_adr = 32'h207b0; force soc.dbg_do = 32'h00700493; #1000;
force soc.dbg_adr = 32'h207b4; force soc.dbg_do = 32'h000247b7; #1000;
force soc.dbg_adr = 32'h207b8; force soc.dbg_do = 32'hd3878593; #1000;
force soc.dbg_adr = 32'h207bc; force soc.dbg_do = 32'h00012783; #1000;
force soc.dbg_adr = 32'h207c0; force soc.dbg_do = 32'h04100713; #1000;
force soc.dbg_adr = 32'h207c4; force soc.dbg_do = 32'h00090513; #1000;
force soc.dbg_adr = 32'h207c8; force soc.dbg_do = 32'hbee78aa3; #1000;
force soc.dbg_adr = 32'h207cc; force soc.dbg_do = 32'h04200793; #1000;
force soc.dbg_adr = 32'h207d0; force soc.dbg_do = 32'hbef98a23; #1000;
force soc.dbg_adr = 32'h207d4; force soc.dbg_do = 32'hbf8aac23; #1000;
force soc.dbg_adr = 32'h207d8; force soc.dbg_do = 32'h6f0000ef; #1000;
force soc.dbg_adr = 32'h207dc; force soc.dbg_do = 32'h01214683; #1000;
force soc.dbg_adr = 32'h207e0; force soc.dbg_do = 32'h03314783; #1000;
force soc.dbg_adr = 32'h207e4; force soc.dbg_do = 32'h0ef68063; #1000;
force soc.dbg_adr = 32'h207e8; force soc.dbg_do = 32'h00090593; #1000;
force soc.dbg_adr = 32'h207ec; force soc.dbg_do = 32'h01010513; #1000;
force soc.dbg_adr = 32'h207f0; force soc.dbg_do = 32'h788000ef; #1000;
force soc.dbg_adr = 32'h207f4; force soc.dbg_do = 32'h65cda683; #1000;
force soc.dbg_adr = 32'h207f8; force soc.dbg_do = 32'h00050613; #1000;
force soc.dbg_adr = 32'h207fc; force soc.dbg_do = 32'hc04b2503; #1000;
force soc.dbg_adr = 32'h20800; force soc.dbg_do = 32'h00800793; #1000;
force soc.dbg_adr = 32'h20804; force soc.dbg_do = 32'h00162613; #1000;
force soc.dbg_adr = 32'h20808; force soc.dbg_do = 32'h00168693; #1000;
force soc.dbg_adr = 32'h2080c; force soc.dbg_do = 32'h00500593; #1000;
force soc.dbg_adr = 32'h20810; force soc.dbg_do = 32'hbecaac23; #1000;
force soc.dbg_adr = 32'h20814; force soc.dbg_do = 32'h64ddae23; #1000;
force soc.dbg_adr = 32'h20818; force soc.dbg_do = 32'hbeba2e23; #1000;
force soc.dbg_adr = 32'h2081c; force soc.dbg_do = 32'h08f42c23; #1000;
force soc.dbg_adr = 32'h20820; force soc.dbg_do = 32'h66fda023; #1000;
force soc.dbg_adr = 32'h20824; force soc.dbg_do = 32'h66fda223; #1000;
force soc.dbg_adr = 32'h20828; force soc.dbg_do = 32'h02942023; #1000;
force soc.dbg_adr = 32'h2082c; force soc.dbg_do = 32'h02942223; #1000;
force soc.dbg_adr = 32'h20830; force soc.dbg_do = 32'h609ba023; #1000;
force soc.dbg_adr = 32'h20834; force soc.dbg_do = 32'hca1ff0ef; #1000;
force soc.dbg_adr = 32'h20838; force soc.dbg_do = 32'hbf49c683; #1000;
force soc.dbg_adr = 32'h2083c; force soc.dbg_do = 32'h04000613; #1000;
force soc.dbg_adr = 32'h20840; force soc.dbg_do = 32'h04100793; #1000;
force soc.dbg_adr = 32'h20844; force soc.dbg_do = 32'h00000593; #1000;
force soc.dbg_adr = 32'h20848; force soc.dbg_do = 32'h08d67063; #1000;
force soc.dbg_adr = 32'h2084c; force soc.dbg_do = 32'h00178613; #1000;
force soc.dbg_adr = 32'h20850; force soc.dbg_do = 32'h03858263; #1000;
force soc.dbg_adr = 32'h20854; force soc.dbg_do = 32'h0ff67793; #1000;
force soc.dbg_adr = 32'h20858; force soc.dbg_do = 32'h3cf6e463; #1000;
force soc.dbg_adr = 32'h2085c; force soc.dbg_do = 32'hff9798e3; #1000;
force soc.dbg_adr = 32'h20860; force soc.dbg_do = 32'h00012703; #1000;
force soc.dbg_adr = 32'h20864; force soc.dbg_do = 32'h00100593; #1000;
force soc.dbg_adr = 32'h20868; force soc.dbg_do = 32'h00178613; #1000;
force soc.dbg_adr = 32'h2086c; force soc.dbg_do = 32'hbef70aa3; #1000;
force soc.dbg_adr = 32'h20870; force soc.dbg_do = 32'hff8592e3; #1000;
force soc.dbg_adr = 32'h20874; force soc.dbg_do = 32'h00f12223; #1000;
force soc.dbg_adr = 32'h20878; force soc.dbg_do = 32'h000247b7; #1000;
force soc.dbg_adr = 32'h2087c; force soc.dbg_do = 32'hd5878593; #1000;
force soc.dbg_adr = 32'h20880; force soc.dbg_do = 32'h00090513; #1000;
force soc.dbg_adr = 32'h20884; force soc.dbg_do = 32'h644000ef; #1000;
force soc.dbg_adr = 32'h20888; force soc.dbg_do = 32'h00412783; #1000;
force soc.dbg_adr = 32'h2088c; force soc.dbg_do = 32'hbf49c683; #1000;
force soc.dbg_adr = 32'h20890; force soc.dbg_do = 32'hbfaa2e23; #1000;
force soc.dbg_adr = 32'h20894; force soc.dbg_do = 32'h00178793; #1000;
force soc.dbg_adr = 32'h20898; force soc.dbg_do = 32'h0ff7f793; #1000;
force soc.dbg_adr = 32'h2089c; force soc.dbg_do = 32'h00f6ee63; #1000;
force soc.dbg_adr = 32'h208a0; force soc.dbg_do = 32'hfd979ae3; #1000;
force soc.dbg_adr = 32'h208a4; force soc.dbg_do = 32'h00012703; #1000;
force soc.dbg_adr = 32'h208a8; force soc.dbg_do = 32'hbef70aa3; #1000;
force soc.dbg_adr = 32'h208ac; force soc.dbg_do = 32'h04300713; #1000;
force soc.dbg_adr = 32'h208b0; force soc.dbg_do = 32'h04400793; #1000;
force soc.dbg_adr = 32'h208b4; force soc.dbg_do = 32'hfcd760e3; #1000;
force soc.dbg_adr = 32'h208b8; force soc.dbg_do = 32'h000d0793; #1000;
force soc.dbg_adr = 32'h208bc; force soc.dbg_do = 32'h00012223; #1000;
force soc.dbg_adr = 32'h208c0; force soc.dbg_do = 32'h36c0006f; #1000;
force soc.dbg_adr = 32'h208c4; force soc.dbg_do = 32'h0000006f; #1000;
force soc.dbg_adr = 32'h208c8; force soc.dbg_do = 32'h00100793; #1000;
force soc.dbg_adr = 32'h208cc; force soc.dbg_do = 32'h00f12223; #1000;
force soc.dbg_adr = 32'h208d0; force soc.dbg_do = 32'h00d00693; #1000;
force soc.dbg_adr = 32'h208d4; force soc.dbg_do = 32'h00012703; #1000;
force soc.dbg_adr = 32'h208d8; force soc.dbg_do = 32'hbf574603; #1000;
force soc.dbg_adr = 32'h208dc; force soc.dbg_do = 32'h04100713; #1000;
force soc.dbg_adr = 32'h208e0; force soc.dbg_do = 32'h00e61863; #1000;
force soc.dbg_adr = 32'h208e4; force soc.dbg_do = 32'hbfca2603; #1000;
force soc.dbg_adr = 32'h208e8; force soc.dbg_do = 32'h00978793; #1000;
force soc.dbg_adr = 32'h208ec; force soc.dbg_do = 32'h40c787b3; #1000;
force soc.dbg_adr = 32'h208f0; force soc.dbg_do = 32'h00c12703; #1000;
force soc.dbg_adr = 32'h208f4; force soc.dbg_do = 32'h001d0d13; #1000;
force soc.dbg_adr = 32'h208f8; force soc.dbg_do = 32'heba75ee3; #1000;
force soc.dbg_adr = 32'h208fc; force soc.dbg_do = 32'h06012d03; #1000;
force soc.dbg_adr = 32'h20900; force soc.dbg_do = 32'h00d12623; #1000;
force soc.dbg_adr = 32'h20904; force soc.dbg_do = 32'h00f12423; #1000;
force soc.dbg_adr = 32'h20908; force soc.dbg_do = 32'h829ff0ef; #1000;
force soc.dbg_adr = 32'h2090c; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20910; force soc.dbg_do = 32'hd7850513; #1000;
force soc.dbg_adr = 32'h20914; force soc.dbg_do = 32'h405010ef; #1000;
force soc.dbg_adr = 32'h20918; force soc.dbg_do = 32'h00024cb7; #1000;
force soc.dbg_adr = 32'h2091c; force soc.dbg_do = 32'hbc4c8513; #1000;
force soc.dbg_adr = 32'h20920; force soc.dbg_do = 32'h3f9010ef; #1000;
force soc.dbg_adr = 32'h20924; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20928; force soc.dbg_do = 32'hd8850513; #1000;
force soc.dbg_adr = 32'h2092c; force soc.dbg_do = 32'h3ed010ef; #1000;
force soc.dbg_adr = 32'h20930; force soc.dbg_do = 32'hbc4c8513; #1000;
force soc.dbg_adr = 32'h20934; force soc.dbg_do = 32'h3e5010ef; #1000;
force soc.dbg_adr = 32'h20938; force soc.dbg_do = 32'hbfca2583; #1000;
force soc.dbg_adr = 32'h2093c; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20940; force soc.dbg_do = 32'hdc050513; #1000;
force soc.dbg_adr = 32'h20944; force soc.dbg_do = 32'h000244b7; #1000;
force soc.dbg_adr = 32'h20948; force soc.dbg_do = 32'h3d1010ef; #1000;
force soc.dbg_adr = 32'h2094c; force soc.dbg_do = 32'hddc48513; #1000;
force soc.dbg_adr = 32'h20950; force soc.dbg_do = 32'h00500593; #1000;
force soc.dbg_adr = 32'h20954; force soc.dbg_do = 32'h3c5010ef; #1000;
force soc.dbg_adr = 32'h20958; force soc.dbg_do = 32'hbf8aa583; #1000;
force soc.dbg_adr = 32'h2095c; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20960; force soc.dbg_do = 32'hdf850513; #1000;
force soc.dbg_adr = 32'h20964; force soc.dbg_do = 32'h3b5010ef; #1000;
force soc.dbg_adr = 32'h20968; force soc.dbg_do = 32'hddc48513; #1000;
force soc.dbg_adr = 32'h2096c; force soc.dbg_do = 32'h00100593; #1000;
force soc.dbg_adr = 32'h20970; force soc.dbg_do = 32'h3a9010ef; #1000;
force soc.dbg_adr = 32'h20974; force soc.dbg_do = 32'h00012783; #1000;
force soc.dbg_adr = 32'h20978; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h2097c; force soc.dbg_do = 32'he1450513; #1000;
force soc.dbg_adr = 32'h20980; force soc.dbg_do = 32'hbf57c583; #1000;
force soc.dbg_adr = 32'h20984; force soc.dbg_do = 32'h00024a37; #1000;
force soc.dbg_adr = 32'h20988; force soc.dbg_do = 32'h00024c37; #1000;
force soc.dbg_adr = 32'h2098c; force soc.dbg_do = 32'h38d010ef; #1000;
force soc.dbg_adr = 32'h20990; force soc.dbg_do = 32'he30a0513; #1000;
force soc.dbg_adr = 32'h20994; force soc.dbg_do = 32'h04100593; #1000;
force soc.dbg_adr = 32'h20998; force soc.dbg_do = 32'h381010ef; #1000;
force soc.dbg_adr = 32'h2099c; force soc.dbg_do = 32'hbf49c583; #1000;
force soc.dbg_adr = 32'h209a0; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h209a4; force soc.dbg_do = 32'he4c50513; #1000;
force soc.dbg_adr = 32'h209a8; force soc.dbg_do = 32'h371010ef; #1000;
force soc.dbg_adr = 32'h209ac; force soc.dbg_do = 32'he30a0513; #1000;
force soc.dbg_adr = 32'h209b0; force soc.dbg_do = 32'h04200593; #1000;
force soc.dbg_adr = 32'h209b4; force soc.dbg_do = 32'h365010ef; #1000;
force soc.dbg_adr = 32'h209b8; force soc.dbg_do = 32'h02042583; #1000;
force soc.dbg_adr = 32'h209bc; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h209c0; force soc.dbg_do = 32'he6850513; #1000;
force soc.dbg_adr = 32'h209c4; force soc.dbg_do = 32'h355010ef; #1000;
force soc.dbg_adr = 32'h209c8; force soc.dbg_do = 32'hddc48513; #1000;
force soc.dbg_adr = 32'h209cc; force soc.dbg_do = 32'h00700593; #1000;
force soc.dbg_adr = 32'h209d0; force soc.dbg_do = 32'h349010ef; #1000;
force soc.dbg_adr = 32'h209d4; force soc.dbg_do = 32'h65cda583; #1000;
force soc.dbg_adr = 32'h209d8; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h209dc; force soc.dbg_do = 32'he8450513; #1000;
force soc.dbg_adr = 32'h209e0; force soc.dbg_do = 32'h339010ef; #1000;
force soc.dbg_adr = 32'h209e4; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h209e8; force soc.dbg_do = 32'hea050513; #1000;
force soc.dbg_adr = 32'h209ec; force soc.dbg_do = 32'h32d010ef; #1000;
force soc.dbg_adr = 32'h209f0; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h209f4; force soc.dbg_do = 32'hecc50513; #1000;
force soc.dbg_adr = 32'h209f8; force soc.dbg_do = 32'h321010ef; #1000;
force soc.dbg_adr = 32'h209fc; force soc.dbg_do = 32'hc04b2703; #1000;
force soc.dbg_adr = 32'h20a00; force soc.dbg_do = 32'hed8c0513; #1000;
force soc.dbg_adr = 32'h20a04; force soc.dbg_do = 32'h00024bb7; #1000;
force soc.dbg_adr = 32'h20a08; force soc.dbg_do = 32'h00072583; #1000;
force soc.dbg_adr = 32'h20a0c; force soc.dbg_do = 32'h00024ab7; #1000;
force soc.dbg_adr = 32'h20a10; force soc.dbg_do = 32'h00024a37; #1000;
force soc.dbg_adr = 32'h20a14; force soc.dbg_do = 32'h305010ef; #1000;
force soc.dbg_adr = 32'h20a18; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20a1c; force soc.dbg_do = 32'hef450513; #1000;
force soc.dbg_adr = 32'h20a20; force soc.dbg_do = 32'h2f9010ef; #1000;
force soc.dbg_adr = 32'h20a24; force soc.dbg_do = 32'hc04b2703; #1000;
force soc.dbg_adr = 32'h20a28; force soc.dbg_do = 32'hf28b8513; #1000;
force soc.dbg_adr = 32'h20a2c; force soc.dbg_do = 32'h000249b7; #1000;
force soc.dbg_adr = 32'h20a30; force soc.dbg_do = 32'h00472583; #1000;
force soc.dbg_adr = 32'h20a34; force soc.dbg_do = 32'h00024437; #1000;
force soc.dbg_adr = 32'h20a38; force soc.dbg_do = 32'h2e1010ef; #1000;
force soc.dbg_adr = 32'h20a3c; force soc.dbg_do = 32'hddc48513; #1000;
force soc.dbg_adr = 32'h20a40; force soc.dbg_do = 32'h00000593; #1000;
force soc.dbg_adr = 32'h20a44; force soc.dbg_do = 32'h2d5010ef; #1000;
force soc.dbg_adr = 32'h20a48; force soc.dbg_do = 32'hc04b2703; #1000;
force soc.dbg_adr = 32'h20a4c; force soc.dbg_do = 32'hf44a8513; #1000;
force soc.dbg_adr = 32'h20a50; force soc.dbg_do = 32'h00872583; #1000;
force soc.dbg_adr = 32'h20a54; force soc.dbg_do = 32'h2c5010ef; #1000;
force soc.dbg_adr = 32'h20a58; force soc.dbg_do = 32'hddc48513; #1000;
force soc.dbg_adr = 32'h20a5c; force soc.dbg_do = 32'h00200593; #1000;
force soc.dbg_adr = 32'h20a60; force soc.dbg_do = 32'h2b9010ef; #1000;
force soc.dbg_adr = 32'h20a64; force soc.dbg_do = 32'hc04b2703; #1000;
force soc.dbg_adr = 32'h20a68; force soc.dbg_do = 32'hf60a0513; #1000;
force soc.dbg_adr = 32'h20a6c; force soc.dbg_do = 32'h00c72583; #1000;
force soc.dbg_adr = 32'h20a70; force soc.dbg_do = 32'h2a9010ef; #1000;
force soc.dbg_adr = 32'h20a74; force soc.dbg_do = 32'hddc48513; #1000;
force soc.dbg_adr = 32'h20a78; force soc.dbg_do = 32'h01100593; #1000;
force soc.dbg_adr = 32'h20a7c; force soc.dbg_do = 32'h29d010ef; #1000;
force soc.dbg_adr = 32'h20a80; force soc.dbg_do = 32'hc04b2583; #1000;
force soc.dbg_adr = 32'h20a84; force soc.dbg_do = 32'hf7c98513; #1000;
force soc.dbg_adr = 32'h20a88; force soc.dbg_do = 32'h00003b37; #1000;
force soc.dbg_adr = 32'h20a8c; force soc.dbg_do = 32'h01058593; #1000;
force soc.dbg_adr = 32'h20a90; force soc.dbg_do = 32'h289010ef; #1000;
force soc.dbg_adr = 32'h20a94; force soc.dbg_do = 32'hf9840513; #1000;
force soc.dbg_adr = 32'h20a98; force soc.dbg_do = 32'h281010ef; #1000;
force soc.dbg_adr = 32'h20a9c; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20aa0; force soc.dbg_do = 32'hfd050513; #1000;
force soc.dbg_adr = 32'h20aa4; force soc.dbg_do = 32'h275010ef; #1000;
force soc.dbg_adr = 32'h20aa8; force soc.dbg_do = 32'hc00b2703; #1000;
force soc.dbg_adr = 32'h20aac; force soc.dbg_do = 32'hed8c0513; #1000;
force soc.dbg_adr = 32'h20ab0; force soc.dbg_do = 32'h00072583; #1000;
force soc.dbg_adr = 32'h20ab4; force soc.dbg_do = 32'h265010ef; #1000;
force soc.dbg_adr = 32'h20ab8; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20abc; force soc.dbg_do = 32'hfe450513; #1000;
force soc.dbg_adr = 32'h20ac0; force soc.dbg_do = 32'h259010ef; #1000;
force soc.dbg_adr = 32'h20ac4; force soc.dbg_do = 32'hc00b2703; #1000;
force soc.dbg_adr = 32'h20ac8; force soc.dbg_do = 32'hf28b8513; #1000;
force soc.dbg_adr = 32'h20acc; force soc.dbg_do = 32'h00472583; #1000;
force soc.dbg_adr = 32'h20ad0; force soc.dbg_do = 32'h249010ef; #1000;
force soc.dbg_adr = 32'h20ad4; force soc.dbg_do = 32'hddc48513; #1000;
force soc.dbg_adr = 32'h20ad8; force soc.dbg_do = 32'h00000593; #1000;
force soc.dbg_adr = 32'h20adc; force soc.dbg_do = 32'h23d010ef; #1000;
force soc.dbg_adr = 32'h20ae0; force soc.dbg_do = 32'hc00b2703; #1000;
force soc.dbg_adr = 32'h20ae4; force soc.dbg_do = 32'hf44a8513; #1000;
force soc.dbg_adr = 32'h20ae8; force soc.dbg_do = 32'h00872583; #1000;
force soc.dbg_adr = 32'h20aec; force soc.dbg_do = 32'h22d010ef; #1000;
force soc.dbg_adr = 32'h20af0; force soc.dbg_do = 32'hddc48513; #1000;
force soc.dbg_adr = 32'h20af4; force soc.dbg_do = 32'h00100593; #1000;
force soc.dbg_adr = 32'h20af8; force soc.dbg_do = 32'h221010ef; #1000;
force soc.dbg_adr = 32'h20afc; force soc.dbg_do = 32'hc00b2703; #1000;
force soc.dbg_adr = 32'h20b00; force soc.dbg_do = 32'hf60a0513; #1000;
force soc.dbg_adr = 32'h20b04; force soc.dbg_do = 32'h00c72583; #1000;
force soc.dbg_adr = 32'h20b08; force soc.dbg_do = 32'h211010ef; #1000;
force soc.dbg_adr = 32'h20b0c; force soc.dbg_do = 32'hddc48513; #1000;
force soc.dbg_adr = 32'h20b10; force soc.dbg_do = 32'h01200593; #1000;
force soc.dbg_adr = 32'h20b14; force soc.dbg_do = 32'h205010ef; #1000;
force soc.dbg_adr = 32'h20b18; force soc.dbg_do = 32'hc00b2583; #1000;
force soc.dbg_adr = 32'h20b1c; force soc.dbg_do = 32'hf7c98513; #1000;
force soc.dbg_adr = 32'h20b20; force soc.dbg_do = 32'h01058593; #1000;
force soc.dbg_adr = 32'h20b24; force soc.dbg_do = 32'h1f5010ef; #1000;
force soc.dbg_adr = 32'h20b28; force soc.dbg_do = 32'hf9840513; #1000;
force soc.dbg_adr = 32'h20b2c; force soc.dbg_do = 32'h1ed010ef; #1000;
force soc.dbg_adr = 32'h20b30; force soc.dbg_do = 32'h00812783; #1000;
force soc.dbg_adr = 32'h20b34; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20b38; force soc.dbg_do = 32'h02450513; #1000;
force soc.dbg_adr = 32'h20b3c; force soc.dbg_do = 32'h00078593; #1000;
force soc.dbg_adr = 32'h20b40; force soc.dbg_do = 32'h1d9010ef; #1000;
force soc.dbg_adr = 32'h20b44; force soc.dbg_do = 32'hddc48513; #1000;
force soc.dbg_adr = 32'h20b48; force soc.dbg_do = 32'h00500593; #1000;
force soc.dbg_adr = 32'h20b4c; force soc.dbg_do = 32'h1cd010ef; #1000;
force soc.dbg_adr = 32'h20b50; force soc.dbg_do = 32'h00c12683; #1000;
force soc.dbg_adr = 32'h20b54; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20b58; force soc.dbg_do = 32'h04050513; #1000;
force soc.dbg_adr = 32'h20b5c; force soc.dbg_do = 32'h00068593; #1000;
force soc.dbg_adr = 32'h20b60; force soc.dbg_do = 32'h1b9010ef; #1000;
force soc.dbg_adr = 32'h20b64; force soc.dbg_do = 32'hddc48513; #1000;
force soc.dbg_adr = 32'h20b68; force soc.dbg_do = 32'h00d00593; #1000;
force soc.dbg_adr = 32'h20b6c; force soc.dbg_do = 32'h1ad010ef; #1000;
force soc.dbg_adr = 32'h20b70; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20b74; force soc.dbg_do = 32'h00700593; #1000;
force soc.dbg_adr = 32'h20b78; force soc.dbg_do = 32'h05c50513; #1000;
force soc.dbg_adr = 32'h20b7c; force soc.dbg_do = 32'h19d010ef; #1000;
force soc.dbg_adr = 32'h20b80; force soc.dbg_do = 32'hddc48513; #1000;
force soc.dbg_adr = 32'h20b84; force soc.dbg_do = 32'h00700593; #1000;
force soc.dbg_adr = 32'h20b88; force soc.dbg_do = 32'h191010ef; #1000;
force soc.dbg_adr = 32'h20b8c; force soc.dbg_do = 32'h00412583; #1000;
force soc.dbg_adr = 32'h20b90; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20b94; force soc.dbg_do = 32'h07850513; #1000;
force soc.dbg_adr = 32'h20b98; force soc.dbg_do = 32'h181010ef; #1000;
force soc.dbg_adr = 32'h20b9c; force soc.dbg_do = 32'hddc48513; #1000;
force soc.dbg_adr = 32'h20ba0; force soc.dbg_do = 32'h00100593; #1000;
force soc.dbg_adr = 32'h20ba4; force soc.dbg_do = 32'h175010ef; #1000;
force soc.dbg_adr = 32'h20ba8; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20bac; force soc.dbg_do = 32'h01010593; #1000;
force soc.dbg_adr = 32'h20bb0; force soc.dbg_do = 32'h09450513; #1000;
force soc.dbg_adr = 32'h20bb4; force soc.dbg_do = 32'h165010ef; #1000;
force soc.dbg_adr = 32'h20bb8; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20bbc; force soc.dbg_do = 32'h0b050513; #1000;
force soc.dbg_adr = 32'h20bc0; force soc.dbg_do = 32'h159010ef; #1000;
force soc.dbg_adr = 32'h20bc4; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20bc8; force soc.dbg_do = 32'h00090593; #1000;
force soc.dbg_adr = 32'h20bcc; force soc.dbg_do = 32'h0e850513; #1000;
force soc.dbg_adr = 32'h20bd0; force soc.dbg_do = 32'h149010ef; #1000;
force soc.dbg_adr = 32'h20bd4; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20bd8; force soc.dbg_do = 32'h10450513; #1000;
force soc.dbg_adr = 32'h20bdc; force soc.dbg_do = 32'h13d010ef; #1000;
force soc.dbg_adr = 32'h20be0; force soc.dbg_do = 32'hbc4c8513; #1000;
force soc.dbg_adr = 32'h20be4; force soc.dbg_do = 32'h135010ef; #1000;
force soc.dbg_adr = 32'h20be8; force soc.dbg_do = 32'h08c12083; #1000;
force soc.dbg_adr = 32'h20bec; force soc.dbg_do = 32'h08812403; #1000;
force soc.dbg_adr = 32'h20bf0; force soc.dbg_do = 32'h08412483; #1000;
force soc.dbg_adr = 32'h20bf4; force soc.dbg_do = 32'h08012903; #1000;
force soc.dbg_adr = 32'h20bf8; force soc.dbg_do = 32'h07c12983; #1000;
force soc.dbg_adr = 32'h20bfc; force soc.dbg_do = 32'h07812a03; #1000;
force soc.dbg_adr = 32'h20c00; force soc.dbg_do = 32'h07412a83; #1000;
force soc.dbg_adr = 32'h20c04; force soc.dbg_do = 32'h07012b03; #1000;
force soc.dbg_adr = 32'h20c08; force soc.dbg_do = 32'h06c12b83; #1000;
force soc.dbg_adr = 32'h20c0c; force soc.dbg_do = 32'h06812c03; #1000;
force soc.dbg_adr = 32'h20c10; force soc.dbg_do = 32'h06412c83; #1000;
force soc.dbg_adr = 32'h20c14; force soc.dbg_do = 32'h05c12d83; #1000;
force soc.dbg_adr = 32'h20c18; force soc.dbg_do = 32'h09010113; #1000;
force soc.dbg_adr = 32'h20c1c; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20c20; force soc.dbg_do = 32'h00100793; #1000;
force soc.dbg_adr = 32'h20c24; force soc.dbg_do = 32'h00f12223; #1000;
force soc.dbg_adr = 32'h20c28; force soc.dbg_do = 32'h00300793; #1000;
force soc.dbg_adr = 32'h20c2c; force soc.dbg_do = 32'h00179693; #1000;
force soc.dbg_adr = 32'h20c30; force soc.dbg_do = 32'h00f686b3; #1000;
force soc.dbg_adr = 32'h20c34; force soc.dbg_do = 32'h00068513; #1000;
force soc.dbg_adr = 32'h20c38; force soc.dbg_do = 32'h00700593; #1000;
force soc.dbg_adr = 32'h20c3c; force soc.dbg_do = 32'h00d12423; #1000;
force soc.dbg_adr = 32'h20c40; force soc.dbg_do = 32'h635020ef; #1000;
force soc.dbg_adr = 32'h20c44; force soc.dbg_do = 32'h00812683; #1000;
force soc.dbg_adr = 32'h20c48; force soc.dbg_do = 32'h00050793; #1000;
force soc.dbg_adr = 32'h20c4c; force soc.dbg_do = 32'hff968693; #1000;
force soc.dbg_adr = 32'h20c50; force soc.dbg_do = 32'h00369613; #1000;
force soc.dbg_adr = 32'h20c54; force soc.dbg_do = 32'h40d606b3; #1000;
force soc.dbg_adr = 32'h20c58; force soc.dbg_do = 32'h40a686b3; #1000;
force soc.dbg_adr = 32'h20c5c; force soc.dbg_do = 32'hc79ff06f; #1000;
force soc.dbg_adr = 32'h20c60; force soc.dbg_do = 32'h00024537; #1000;
force soc.dbg_adr = 32'h20c64; force soc.dbg_do = 32'hcd850513; #1000;
force soc.dbg_adr = 32'h20c68; force soc.dbg_do = 32'h00d12423; #1000;
force soc.dbg_adr = 32'h20c6c; force soc.dbg_do = 32'h00f12023; #1000;
force soc.dbg_adr = 32'h20c70; force soc.dbg_do = 32'h0a9010ef; #1000;
force soc.dbg_adr = 32'h20c74; force soc.dbg_do = 32'h000247b7; #1000;
force soc.dbg_adr = 32'h20c78; force soc.dbg_do = 32'hbc478513; #1000;
force soc.dbg_adr = 32'h20c7c; force soc.dbg_do = 32'h09d010ef; #1000;
force soc.dbg_adr = 32'h20c80; force soc.dbg_do = 32'h00812683; #1000;
force soc.dbg_adr = 32'h20c84; force soc.dbg_do = 32'h00012783; #1000;
force soc.dbg_adr = 32'h20c88; force soc.dbg_do = 32'hac9ff06f; #1000;
force soc.dbg_adr = 32'h20c8c; force soc.dbg_do = 32'h00003737; #1000;
force soc.dbg_adr = 32'h20c90; force soc.dbg_do = 32'h00000413; #1000;
force soc.dbg_adr = 32'h20c94; force soc.dbg_do = 32'h00e12023; #1000;
force soc.dbg_adr = 32'h20c98; force soc.dbg_do = 32'h00003ab7; #1000;
force soc.dbg_adr = 32'h20c9c; force soc.dbg_do = 32'h000039b7; #1000;
force soc.dbg_adr = 32'h20ca0; force soc.dbg_do = 32'h03010913; #1000;
force soc.dbg_adr = 32'h20ca4; force soc.dbg_do = 32'h00003a37; #1000;
force soc.dbg_adr = 32'h20ca8; force soc.dbg_do = 32'hc59ff06f; #1000;
force soc.dbg_adr = 32'h20cac; force soc.dbg_do = 32'h000037b7; #1000;
force soc.dbg_adr = 32'h20cb0; force soc.dbg_do = 32'hbf57c703; #1000;
force soc.dbg_adr = 32'h20cb4; force soc.dbg_do = 32'h04100793; #1000;
force soc.dbg_adr = 32'h20cb8; force soc.dbg_do = 32'h00f70463; #1000;
force soc.dbg_adr = 32'h20cbc; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20cc0; force soc.dbg_do = 32'h00052783; #1000;
force soc.dbg_adr = 32'h20cc4; force soc.dbg_do = 32'h00003737; #1000;
force soc.dbg_adr = 32'h20cc8; force soc.dbg_do = 32'hbfc72703; #1000;
force soc.dbg_adr = 32'h20ccc; force soc.dbg_do = 32'h00978793; #1000;
force soc.dbg_adr = 32'h20cd0; force soc.dbg_do = 32'h40e787b3; #1000;
force soc.dbg_adr = 32'h20cd4; force soc.dbg_do = 32'h00f52023; #1000;
force soc.dbg_adr = 32'h20cd8; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20cdc; force soc.dbg_do = 32'h00003737; #1000;
force soc.dbg_adr = 32'h20ce0; force soc.dbg_do = 32'hc0472783; #1000;
force soc.dbg_adr = 32'h20ce4; force soc.dbg_do = 32'h00078863; #1000;
force soc.dbg_adr = 32'h20ce8; force soc.dbg_do = 32'h0007a783; #1000;
force soc.dbg_adr = 32'h20cec; force soc.dbg_do = 32'h00f52023; #1000;
force soc.dbg_adr = 32'h20cf0; force soc.dbg_do = 32'hc0472783; #1000;
force soc.dbg_adr = 32'h20cf4; force soc.dbg_do = 32'h00003737; #1000;
force soc.dbg_adr = 32'h20cf8; force soc.dbg_do = 32'hbfc72703; #1000;
force soc.dbg_adr = 32'h20cfc; force soc.dbg_do = 32'h00c70713; #1000;
force soc.dbg_adr = 32'h20d00; force soc.dbg_do = 32'h00e7a623; #1000;
force soc.dbg_adr = 32'h20d04; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20d08; force soc.dbg_do = 32'h000037b7; #1000;
force soc.dbg_adr = 32'h20d0c; force soc.dbg_do = 32'hbf57c783; #1000;
force soc.dbg_adr = 32'h20d10; force soc.dbg_do = 32'h00003737; #1000;
force soc.dbg_adr = 32'h20d14; force soc.dbg_do = 32'hbf872683; #1000;
force soc.dbg_adr = 32'h20d18; force soc.dbg_do = 32'hfbf78793; #1000;
force soc.dbg_adr = 32'h20d1c; force soc.dbg_do = 32'h0017b793; #1000;
force soc.dbg_adr = 32'h20d20; force soc.dbg_do = 32'h00d7e7b3; #1000;
force soc.dbg_adr = 32'h20d24; force soc.dbg_do = 32'h04200613; #1000;
force soc.dbg_adr = 32'h20d28; force soc.dbg_do = 32'h000036b7; #1000;
force soc.dbg_adr = 32'h20d2c; force soc.dbg_do = 32'hbef72c23; #1000;
force soc.dbg_adr = 32'h20d30; force soc.dbg_do = 32'hbec68a23; #1000;
force soc.dbg_adr = 32'h20d34; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20d38; force soc.dbg_do = 32'h00003737; #1000;
force soc.dbg_adr = 32'h20d3c; force soc.dbg_do = 32'h04100693; #1000;
force soc.dbg_adr = 32'h20d40; force soc.dbg_do = 32'h000037b7; #1000;
force soc.dbg_adr = 32'h20d44; force soc.dbg_do = 32'hbed70aa3; #1000;
force soc.dbg_adr = 32'h20d48; force soc.dbg_do = 32'hbe07ac23; #1000;
force soc.dbg_adr = 32'h20d4c; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20d50; force soc.dbg_do = 32'h00200793; #1000;
force soc.dbg_adr = 32'h20d54; force soc.dbg_do = 32'h02f50e63; #1000;
force soc.dbg_adr = 32'h20d58; force soc.dbg_do = 32'h00300713; #1000;
force soc.dbg_adr = 32'h20d5c; force soc.dbg_do = 32'h00e5a023; #1000;
force soc.dbg_adr = 32'h20d60; force soc.dbg_do = 32'h00100713; #1000;
force soc.dbg_adr = 32'h20d64; force soc.dbg_do = 32'h00e50a63; #1000;
force soc.dbg_adr = 32'h20d68; force soc.dbg_do = 32'h00400713; #1000;
force soc.dbg_adr = 32'h20d6c; force soc.dbg_do = 32'h02e50863; #1000;
force soc.dbg_adr = 32'h20d70; force soc.dbg_do = 32'h00050c63; #1000;
force soc.dbg_adr = 32'h20d74; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20d78; force soc.dbg_do = 32'h000037b7; #1000;
force soc.dbg_adr = 32'h20d7c; force soc.dbg_do = 32'hbfc7a703; #1000;
force soc.dbg_adr = 32'h20d80; force soc.dbg_do = 32'h06400793; #1000;
force soc.dbg_adr = 32'h20d84; force soc.dbg_do = 32'hfee7d8e3; #1000;
force soc.dbg_adr = 32'h20d88; force soc.dbg_do = 32'h0005a023; #1000;
force soc.dbg_adr = 32'h20d8c; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20d90; force soc.dbg_do = 32'h00100793; #1000;
force soc.dbg_adr = 32'h20d94; force soc.dbg_do = 32'h00f5a023; #1000;
force soc.dbg_adr = 32'h20d98; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20d9c; force soc.dbg_do = 32'h00f5a023; #1000;
force soc.dbg_adr = 32'h20da0; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20da4; force soc.dbg_do = 32'h00250513; #1000;
force soc.dbg_adr = 32'h20da8; force soc.dbg_do = 32'h00b50533; #1000;
force soc.dbg_adr = 32'h20dac; force soc.dbg_do = 32'h00a62023; #1000;
force soc.dbg_adr = 32'h20db0; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20db4; force soc.dbg_do = 32'h00560713; #1000;
force soc.dbg_adr = 32'h20db8; force soc.dbg_do = 32'h00171793; #1000;
force soc.dbg_adr = 32'h20dbc; force soc.dbg_do = 32'h00e787b3; #1000;
force soc.dbg_adr = 32'h20dc0; force soc.dbg_do = 32'h00379793; #1000;
force soc.dbg_adr = 32'h20dc4; force soc.dbg_do = 32'h00e787b3; #1000;
force soc.dbg_adr = 32'h20dc8; force soc.dbg_do = 32'h00261613; #1000;
force soc.dbg_adr = 32'h20dcc; force soc.dbg_do = 32'h00271813; #1000;
force soc.dbg_adr = 32'h20dd0; force soc.dbg_do = 32'h00379793; #1000;
force soc.dbg_adr = 32'h20dd4; force soc.dbg_do = 32'h01050533; #1000;
force soc.dbg_adr = 32'h20dd8; force soc.dbg_do = 32'h00f60833; #1000;
force soc.dbg_adr = 32'h20ddc; force soc.dbg_do = 32'h00d52023; #1000;
force soc.dbg_adr = 32'h20de0; force soc.dbg_do = 32'h00d52223; #1000;
force soc.dbg_adr = 32'h20de4; force soc.dbg_do = 32'h06e52c23; #1000;
force soc.dbg_adr = 32'h20de8; force soc.dbg_do = 32'h010586b3; #1000;
force soc.dbg_adr = 32'h20dec; force soc.dbg_do = 32'h0106a803; #1000;
force soc.dbg_adr = 32'h20df0; force soc.dbg_do = 32'h00e6aa23; #1000;
force soc.dbg_adr = 32'h20df4; force soc.dbg_do = 32'h00e6ac23; #1000;
force soc.dbg_adr = 32'h20df8; force soc.dbg_do = 32'h00180713; #1000;
force soc.dbg_adr = 32'h20dfc; force soc.dbg_do = 32'h00e6a823; #1000;
force soc.dbg_adr = 32'h20e00; force soc.dbg_do = 32'h00c585b3; #1000;
force soc.dbg_adr = 32'h20e04; force soc.dbg_do = 32'h00052603; #1000;
force soc.dbg_adr = 32'h20e08; force soc.dbg_do = 32'h00f585b3; #1000;
force soc.dbg_adr = 32'h20e0c; force soc.dbg_do = 32'h000017b7; #1000;
force soc.dbg_adr = 32'h20e10; force soc.dbg_do = 32'h00b787b3; #1000;
force soc.dbg_adr = 32'h20e14; force soc.dbg_do = 32'h00003737; #1000;
force soc.dbg_adr = 32'h20e18; force soc.dbg_do = 32'h00500693; #1000;
force soc.dbg_adr = 32'h20e1c; force soc.dbg_do = 32'hfac7aa23; #1000;
force soc.dbg_adr = 32'h20e20; force soc.dbg_do = 32'hbed72e23; #1000;
force soc.dbg_adr = 32'h20e24; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20e28; force soc.dbg_do = 32'h0ff57513; #1000;
force soc.dbg_adr = 32'h20e2c; force soc.dbg_do = 32'h0ff5f593; #1000;
force soc.dbg_adr = 32'h20e30; force soc.dbg_do = 32'h00b50663; #1000;
force soc.dbg_adr = 32'h20e34; force soc.dbg_do = 32'h00000513; #1000;
force soc.dbg_adr = 32'h20e38; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20e3c; force soc.dbg_do = 32'h000037b7; #1000;
force soc.dbg_adr = 32'h20e40; force soc.dbg_do = 32'hbea78aa3; #1000;
force soc.dbg_adr = 32'h20e44; force soc.dbg_do = 32'h00100513; #1000;
force soc.dbg_adr = 32'h20e48; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20e4c; force soc.dbg_do = 32'h00254703; #1000;
force soc.dbg_adr = 32'h20e50; force soc.dbg_do = 32'h0035c783; #1000;
force soc.dbg_adr = 32'h20e54; force soc.dbg_do = 32'h02f70c63; #1000;
force soc.dbg_adr = 32'h20e58; force soc.dbg_do = 32'hff010113; #1000;
force soc.dbg_adr = 32'h20e5c; force soc.dbg_do = 32'h00112623; #1000;
force soc.dbg_adr = 32'h20e60; force soc.dbg_do = 32'h118000ef; #1000;
force soc.dbg_adr = 32'h20e64; force soc.dbg_do = 32'h00000793; #1000;
force soc.dbg_adr = 32'h20e68; force soc.dbg_do = 32'h00a05a63; #1000;
force soc.dbg_adr = 32'h20e6c; force soc.dbg_do = 32'h000037b7; #1000;
force soc.dbg_adr = 32'h20e70; force soc.dbg_do = 32'h00a00713; #1000;
force soc.dbg_adr = 32'h20e74; force soc.dbg_do = 32'hbee7ae23; #1000;
force soc.dbg_adr = 32'h20e78; force soc.dbg_do = 32'h00100793; #1000;
force soc.dbg_adr = 32'h20e7c; force soc.dbg_do = 32'h00c12083; #1000;
force soc.dbg_adr = 32'h20e80; force soc.dbg_do = 32'h00078513; #1000;
force soc.dbg_adr = 32'h20e84; force soc.dbg_do = 32'h01010113; #1000;
force soc.dbg_adr = 32'h20e88; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20e8c; force soc.dbg_do = 32'h0000006f; #1000;
force soc.dbg_adr = 32'h20e90; force soc.dbg_do = 32'hffe50513; #1000;
force soc.dbg_adr = 32'h20e94; force soc.dbg_do = 32'h00153513; #1000;
force soc.dbg_adr = 32'h20e98; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20e9c; force soc.dbg_do = 32'h00003637; #1000;
force soc.dbg_adr = 32'h20ea0; force soc.dbg_do = 32'hc0862683; #1000;
force soc.dbg_adr = 32'h20ea4; force soc.dbg_do = 32'h000027b7; #1000;
force soc.dbg_adr = 32'h20ea8; force soc.dbg_do = 32'h7d878793; #1000;
force soc.dbg_adr = 32'h20eac; force soc.dbg_do = 32'h00a68733; #1000;
force soc.dbg_adr = 32'h20eb0; force soc.dbg_do = 32'hc0e62423; #1000;
force soc.dbg_adr = 32'h20eb4; force soc.dbg_do = 32'h40000613; #1000;
force soc.dbg_adr = 32'h20eb8; force soc.dbg_do = 32'h00d78533; #1000;
force soc.dbg_adr = 32'h20ebc; force soc.dbg_do = 32'h00e65463; #1000;
force soc.dbg_adr = 32'h20ec0; force soc.dbg_do = 32'h00100073; #1000;
force soc.dbg_adr = 32'h20ec4; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20ec8; force soc.dbg_do = 32'h00050793; #1000;
force soc.dbg_adr = 32'h20ecc; force soc.dbg_do = 32'h0180006f; #1000;
force soc.dbg_adr = 32'h20ed0; force soc.dbg_do = 32'h0005c703; #1000;
force soc.dbg_adr = 32'h20ed4; force soc.dbg_do = 32'h00158593; #1000;
force soc.dbg_adr = 32'h20ed8; force soc.dbg_do = 32'h00178793; #1000;
force soc.dbg_adr = 32'h20edc; force soc.dbg_do = 32'hfee78fa3; #1000;
force soc.dbg_adr = 32'h20ee0; force soc.dbg_do = 32'h08070463; #1000;
force soc.dbg_adr = 32'h20ee4; force soc.dbg_do = 32'h00f5e733; #1000;
force soc.dbg_adr = 32'h20ee8; force soc.dbg_do = 32'h00377713; #1000;
force soc.dbg_adr = 32'h20eec; force soc.dbg_do = 32'hfe0712e3; #1000;
force soc.dbg_adr = 32'h20ef0; force soc.dbg_do = 32'h0005a683; #1000;
force soc.dbg_adr = 32'h20ef4; force soc.dbg_do = 32'hfeff08b7; #1000;
force soc.dbg_adr = 32'h20ef8; force soc.dbg_do = 32'heff88893; #1000;
force soc.dbg_adr = 32'h20efc; force soc.dbg_do = 32'h01168733; #1000;
force soc.dbg_adr = 32'h20f00; force soc.dbg_do = 32'hfff6c613; #1000;
force soc.dbg_adr = 32'h20f04; force soc.dbg_do = 32'h80808837; #1000;
force soc.dbg_adr = 32'h20f08; force soc.dbg_do = 32'h00c77733; #1000;
force soc.dbg_adr = 32'h20f0c; force soc.dbg_do = 32'h08080813; #1000;
force soc.dbg_adr = 32'h20f10; force soc.dbg_do = 32'h01077733; #1000;
force soc.dbg_adr = 32'h20f14; force soc.dbg_do = 32'h02071463; #1000;
force soc.dbg_adr = 32'h20f18; force soc.dbg_do = 32'h00d7a023; #1000;
force soc.dbg_adr = 32'h20f1c; force soc.dbg_do = 32'h0045a683; #1000;
force soc.dbg_adr = 32'h20f20; force soc.dbg_do = 32'h00458593; #1000;
force soc.dbg_adr = 32'h20f24; force soc.dbg_do = 32'h00478793; #1000;
force soc.dbg_adr = 32'h20f28; force soc.dbg_do = 32'h01168733; #1000;
force soc.dbg_adr = 32'h20f2c; force soc.dbg_do = 32'hfff6c613; #1000;
force soc.dbg_adr = 32'h20f30; force soc.dbg_do = 32'h00c77733; #1000;
force soc.dbg_adr = 32'h20f34; force soc.dbg_do = 32'h01077733; #1000;
force soc.dbg_adr = 32'h20f38; force soc.dbg_do = 32'hfe0700e3; #1000;
force soc.dbg_adr = 32'h20f3c; force soc.dbg_do = 32'h00d78023; #1000;
force soc.dbg_adr = 32'h20f40; force soc.dbg_do = 32'h0ff6f713; #1000;
force soc.dbg_adr = 32'h20f44; force soc.dbg_do = 32'h02070263; #1000;
force soc.dbg_adr = 32'h20f48; force soc.dbg_do = 32'h0086d713; #1000;
force soc.dbg_adr = 32'h20f4c; force soc.dbg_do = 32'h00e780a3; #1000;
force soc.dbg_adr = 32'h20f50; force soc.dbg_do = 32'h0ff77713; #1000;
force soc.dbg_adr = 32'h20f54; force soc.dbg_do = 32'h00070a63; #1000;
force soc.dbg_adr = 32'h20f58; force soc.dbg_do = 32'h0106d713; #1000;
force soc.dbg_adr = 32'h20f5c; force soc.dbg_do = 32'h00e78123; #1000;
force soc.dbg_adr = 32'h20f60; force soc.dbg_do = 32'h0ff77713; #1000;
force soc.dbg_adr = 32'h20f64; force soc.dbg_do = 32'h00071463; #1000;
force soc.dbg_adr = 32'h20f68; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20f6c; force soc.dbg_do = 32'h0186d693; #1000;
force soc.dbg_adr = 32'h20f70; force soc.dbg_do = 32'h00d781a3; #1000;
force soc.dbg_adr = 32'h20f74; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20f78; force soc.dbg_do = 32'h01c0006f; #1000;
force soc.dbg_adr = 32'h20f7c; force soc.dbg_do = 32'h00054783; #1000;
force soc.dbg_adr = 32'h20f80; force soc.dbg_do = 32'h0005c703; #1000;
force soc.dbg_adr = 32'h20f84; force soc.dbg_do = 32'h00150513; #1000;
force soc.dbg_adr = 32'h20f88; force soc.dbg_do = 32'h00158593; #1000;
force soc.dbg_adr = 32'h20f8c; force soc.dbg_do = 32'h06e79263; #1000;
force soc.dbg_adr = 32'h20f90; force soc.dbg_do = 32'h04078c63; #1000;
force soc.dbg_adr = 32'h20f94; force soc.dbg_do = 32'h00b567b3; #1000;
force soc.dbg_adr = 32'h20f98; force soc.dbg_do = 32'h0037f793; #1000;
force soc.dbg_adr = 32'h20f9c; force soc.dbg_do = 32'hfe0790e3; #1000;
force soc.dbg_adr = 32'h20fa0; force soc.dbg_do = 32'h00052783; #1000;
force soc.dbg_adr = 32'h20fa4; force soc.dbg_do = 32'h0005a703; #1000;
force soc.dbg_adr = 32'h20fa8; force soc.dbg_do = 32'hfeff0637; #1000;
force soc.dbg_adr = 32'h20fac; force soc.dbg_do = 32'h808086b7; #1000;
force soc.dbg_adr = 32'h20fb0; force soc.dbg_do = 32'heff60613; #1000;
force soc.dbg_adr = 32'h20fb4; force soc.dbg_do = 32'h08068693; #1000;
force soc.dbg_adr = 32'h20fb8; force soc.dbg_do = 32'h00f70a63; #1000;
force soc.dbg_adr = 32'h20fbc; force soc.dbg_do = 32'h0440006f; #1000;
force soc.dbg_adr = 32'h20fc0; force soc.dbg_do = 32'h00052783; #1000;
force soc.dbg_adr = 32'h20fc4; force soc.dbg_do = 32'h0005a703; #1000;
force soc.dbg_adr = 32'h20fc8; force soc.dbg_do = 32'h02e79c63; #1000;
force soc.dbg_adr = 32'h20fcc; force soc.dbg_do = 32'h00c78733; #1000;
force soc.dbg_adr = 32'h20fd0; force soc.dbg_do = 32'hfff7c793; #1000;
force soc.dbg_adr = 32'h20fd4; force soc.dbg_do = 32'h00f777b3; #1000;
force soc.dbg_adr = 32'h20fd8; force soc.dbg_do = 32'h00d7f7b3; #1000;
force soc.dbg_adr = 32'h20fdc; force soc.dbg_do = 32'h00450513; #1000;
force soc.dbg_adr = 32'h20fe0; force soc.dbg_do = 32'h00458593; #1000;
force soc.dbg_adr = 32'h20fe4; force soc.dbg_do = 32'hfc078ee3; #1000;
force soc.dbg_adr = 32'h20fe8; force soc.dbg_do = 32'h00000513; #1000;
force soc.dbg_adr = 32'h20fec; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h20ff0; force soc.dbg_do = 32'h00e7b533; #1000;
force soc.dbg_adr = 32'h20ff4; force soc.dbg_do = 32'h40a00533; #1000;
force soc.dbg_adr = 32'h20ff8; force soc.dbg_do = 32'h00156513; #1000;
force soc.dbg_adr = 32'h20ffc; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h21000; force soc.dbg_do = 32'h0ff7f693; #1000;
force soc.dbg_adr = 32'h21004; force soc.dbg_do = 32'h0ff77613; #1000;
force soc.dbg_adr = 32'h21008; force soc.dbg_do = 32'h04c69c63; #1000;
force soc.dbg_adr = 32'h2100c; force soc.dbg_do = 32'h00000513; #1000;
force soc.dbg_adr = 32'h21010; force soc.dbg_do = 32'hfc068ee3; #1000;
force soc.dbg_adr = 32'h21014; force soc.dbg_do = 32'h0087d693; #1000;
force soc.dbg_adr = 32'h21018; force soc.dbg_do = 32'h00875613; #1000;
force soc.dbg_adr = 32'h2101c; force soc.dbg_do = 32'h0ff6f693; #1000;
force soc.dbg_adr = 32'h21020; force soc.dbg_do = 32'h0ff67613; #1000;
force soc.dbg_adr = 32'h21024; force soc.dbg_do = 32'h02c69e63; #1000;
force soc.dbg_adr = 32'h21028; force soc.dbg_do = 32'hfc0682e3; #1000;
force soc.dbg_adr = 32'h2102c; force soc.dbg_do = 32'h0107d693; #1000;
force soc.dbg_adr = 32'h21030; force soc.dbg_do = 32'h01075613; #1000;
force soc.dbg_adr = 32'h21034; force soc.dbg_do = 32'h0ff6f693; #1000;
force soc.dbg_adr = 32'h21038; force soc.dbg_do = 32'h0ff67613; #1000;
force soc.dbg_adr = 32'h2103c; force soc.dbg_do = 32'h02c69263; #1000;
force soc.dbg_adr = 32'h21040; force soc.dbg_do = 32'hfa0686e3; #1000;
force soc.dbg_adr = 32'h21044; force soc.dbg_do = 32'h0187d793; #1000;
force soc.dbg_adr = 32'h21048; force soc.dbg_do = 32'h01875713; #1000;
force soc.dbg_adr = 32'h2104c; force soc.dbg_do = 32'hfae780e3; #1000;
force soc.dbg_adr = 32'h21050; force soc.dbg_do = 32'h00e7b7b3; #1000;
force soc.dbg_adr = 32'h21054; force soc.dbg_do = 32'h40f007b3; #1000;
force soc.dbg_adr = 32'h21058; force soc.dbg_do = 32'h0017e513; #1000;
force soc.dbg_adr = 32'h2105c; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h21060; force soc.dbg_do = 32'h00c6b7b3; #1000;
force soc.dbg_adr = 32'h21064; force soc.dbg_do = 32'h40f007b3; #1000;
force soc.dbg_adr = 32'h21068; force soc.dbg_do = 32'h0017e513; #1000;
force soc.dbg_adr = 32'h2106c; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h21070; force soc.dbg_do = 32'h00d67663; #1000;
force soc.dbg_adr = 32'h21074; force soc.dbg_do = 32'h00c585b3; #1000;
force soc.dbg_adr = 32'h21078; force soc.dbg_do = 32'h00a58023; #1000;
force soc.dbg_adr = 32'h2107c; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h21080; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h21084; force soc.dbg_do = 32'hfd010113; #1000;
force soc.dbg_adr = 32'h21088; force soc.dbg_do = 32'h03812303; #1000;
force soc.dbg_adr = 32'h2108c; force soc.dbg_do = 32'h02812423; #1000;
force soc.dbg_adr = 32'h21090; force soc.dbg_do = 32'h02912223; #1000;
force soc.dbg_adr = 32'h21094; force soc.dbg_do = 32'h01312e23; #1000;
force soc.dbg_adr = 32'h21098; force soc.dbg_do = 32'h01412c23; #1000;
force soc.dbg_adr = 32'h2109c; force soc.dbg_do = 32'h01512a23; #1000;
force soc.dbg_adr = 32'h210a0; force soc.dbg_do = 32'h01612823; #1000;
force soc.dbg_adr = 32'h210a4; force soc.dbg_do = 32'h01712623; #1000;
force soc.dbg_adr = 32'h210a8; force soc.dbg_do = 32'h01912223; #1000;
force soc.dbg_adr = 32'h210ac; force soc.dbg_do = 32'h02112623; #1000;
force soc.dbg_adr = 32'h210b0; force soc.dbg_do = 32'h03212023; #1000;
force soc.dbg_adr = 32'h210b4; force soc.dbg_do = 32'h01812423; #1000;
force soc.dbg_adr = 32'h210b8; force soc.dbg_do = 32'h00237c93; #1000;
force soc.dbg_adr = 32'h210bc; force soc.dbg_do = 32'h00058a13; #1000;
force soc.dbg_adr = 32'h210c0; force soc.dbg_do = 32'h00070493; #1000;
force soc.dbg_adr = 32'h210c4; force soc.dbg_do = 32'h03412b83; #1000;
force soc.dbg_adr = 32'h210c8; force soc.dbg_do = 32'h03012703; #1000;
force soc.dbg_adr = 32'h210cc; force soc.dbg_do = 32'h00050993; #1000;
force soc.dbg_adr = 32'h210d0; force soc.dbg_do = 32'h00060b13; #1000;
force soc.dbg_adr = 32'h210d4; force soc.dbg_do = 32'h00068a93; #1000;
force soc.dbg_adr = 32'h210d8; force soc.dbg_do = 32'h00078413; #1000;
force soc.dbg_adr = 32'h210dc; force soc.dbg_do = 32'h01037593; #1000;
force soc.dbg_adr = 32'h210e0; force soc.dbg_do = 32'h0e0c8663; #1000;
force soc.dbg_adr = 32'h210e4; force soc.dbg_do = 32'h1c058663; #1000;
force soc.dbg_adr = 32'h210e8; force soc.dbg_do = 32'h40037793; #1000;
force soc.dbg_adr = 32'h210ec; force soc.dbg_do = 32'h1e079e63; #1000;
force soc.dbg_adr = 32'h210f0; force soc.dbg_do = 32'h28041663; #1000;
force soc.dbg_adr = 32'h210f4; force soc.dbg_do = 32'h01000793; #1000;
force soc.dbg_adr = 32'h210f8; force soc.dbg_do = 32'h40f88a63; #1000;
force soc.dbg_adr = 32'h210fc; force soc.dbg_do = 32'h00200793; #1000;
force soc.dbg_adr = 32'h21100; force soc.dbg_do = 32'h42f88863; #1000;
force soc.dbg_adr = 32'h21104; force soc.dbg_do = 32'h03000793; #1000;
force soc.dbg_adr = 32'h21108; force soc.dbg_do = 32'h00f48023; #1000;
force soc.dbg_adr = 32'h2110c; force soc.dbg_do = 32'h00100713; #1000;
force soc.dbg_adr = 32'h21110; force soc.dbg_do = 32'h00337793; #1000;
force soc.dbg_adr = 32'h21114; force soc.dbg_do = 32'h20080e63; #1000;
force soc.dbg_adr = 32'h21118; force soc.dbg_do = 32'h00e486b3; #1000;
force soc.dbg_adr = 32'h2111c; force soc.dbg_do = 32'h02d00613; #1000;
force soc.dbg_adr = 32'h21120; force soc.dbg_do = 32'h00c68023; #1000;
force soc.dbg_adr = 32'h21124; force soc.dbg_do = 32'h00170413; #1000;
force soc.dbg_adr = 32'h21128; force soc.dbg_do = 32'h3c079263; #1000;
force soc.dbg_adr = 32'h2112c; force soc.dbg_do = 32'h11746663; #1000;
force soc.dbg_adr = 32'h21130; force soc.dbg_do = 32'h01a12023; #1000;
force soc.dbg_adr = 32'h21134; force soc.dbg_do = 32'h000b0c13; #1000;
force soc.dbg_adr = 32'h21138; force soc.dbg_do = 32'h008c0c33; #1000;
force soc.dbg_adr = 32'h2113c; force soc.dbg_do = 32'h01848d33; #1000;
force soc.dbg_adr = 32'h21140; force soc.dbg_do = 32'h00848433; #1000;
force soc.dbg_adr = 32'h21144; force soc.dbg_do = 32'hfff44503; #1000;
force soc.dbg_adr = 32'h21148; force soc.dbg_do = 32'h408d0633; #1000;
force soc.dbg_adr = 32'h2114c; force soc.dbg_do = 32'h000a8693; #1000;
force soc.dbg_adr = 32'h21150; force soc.dbg_do = 32'h000a0593; #1000;
force soc.dbg_adr = 32'h21154; force soc.dbg_do = 32'hfff40413; #1000;
force soc.dbg_adr = 32'h21158; force soc.dbg_do = 32'h000c0913; #1000;
force soc.dbg_adr = 32'h2115c; force soc.dbg_do = 32'h000980e7; #1000;
force soc.dbg_adr = 32'h21160; force soc.dbg_do = 32'hfe8492e3; #1000;
force soc.dbg_adr = 32'h21164; force soc.dbg_do = 32'h00012d03; #1000;
force soc.dbg_adr = 32'h21168; force soc.dbg_do = 32'h020c8663; #1000;
force soc.dbg_adr = 32'h2116c; force soc.dbg_do = 32'h41690b33; #1000;
force soc.dbg_adr = 32'h21170; force soc.dbg_do = 32'h037b7263; #1000;
force soc.dbg_adr = 32'h21174; force soc.dbg_do = 32'h00090613; #1000;
force soc.dbg_adr = 32'h21178; force soc.dbg_do = 32'h000a8693; #1000;
force soc.dbg_adr = 32'h2117c; force soc.dbg_do = 32'h000a0593; #1000;
force soc.dbg_adr = 32'h21180; force soc.dbg_do = 32'h02000513; #1000;
force soc.dbg_adr = 32'h21184; force soc.dbg_do = 32'h001b0b13; #1000;
force soc.dbg_adr = 32'h21188; force soc.dbg_do = 32'h00190913; #1000;
force soc.dbg_adr = 32'h2118c; force soc.dbg_do = 32'h000980e7; #1000;
force soc.dbg_adr = 32'h21190; force soc.dbg_do = 32'hff7b62e3; #1000;
force soc.dbg_adr = 32'h21194; force soc.dbg_do = 32'h02c12083; #1000;
force soc.dbg_adr = 32'h21198; force soc.dbg_do = 32'h02812403; #1000;
force soc.dbg_adr = 32'h2119c; force soc.dbg_do = 32'h02412483; #1000;
force soc.dbg_adr = 32'h211a0; force soc.dbg_do = 32'h01c12983; #1000;
force soc.dbg_adr = 32'h211a4; force soc.dbg_do = 32'h01812a03; #1000;
force soc.dbg_adr = 32'h211a8; force soc.dbg_do = 32'h01412a83; #1000;
force soc.dbg_adr = 32'h211ac; force soc.dbg_do = 32'h01012b03; #1000;
force soc.dbg_adr = 32'h211b0; force soc.dbg_do = 32'h00c12b83; #1000;
force soc.dbg_adr = 32'h211b4; force soc.dbg_do = 32'h00812c03; #1000;
force soc.dbg_adr = 32'h211b8; force soc.dbg_do = 32'h00412c83; #1000;
force soc.dbg_adr = 32'h211bc; force soc.dbg_do = 32'h00090513; #1000;
force soc.dbg_adr = 32'h211c0; force soc.dbg_do = 32'h02012903; #1000;
force soc.dbg_adr = 32'h211c4; force soc.dbg_do = 32'h03010113; #1000;
force soc.dbg_adr = 32'h211c8; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h211cc; force soc.dbg_do = 32'h00137513; #1000;
force soc.dbg_adr = 32'h211d0; force soc.dbg_do = 32'h0a0b9c63; #1000;
force soc.dbg_adr = 32'h211d4; force soc.dbg_do = 32'h38e7f263; #1000;
force soc.dbg_adr = 32'h211d8; force soc.dbg_do = 32'h02000693; #1000;
force soc.dbg_adr = 32'h211dc; force soc.dbg_do = 32'h03000613; #1000;
force soc.dbg_adr = 32'h211e0; force soc.dbg_do = 32'h00d40a63; #1000;
force soc.dbg_adr = 32'h211e4; force soc.dbg_do = 32'h00140413; #1000;
force soc.dbg_adr = 32'h211e8; force soc.dbg_do = 32'h008487b3; #1000;
force soc.dbg_adr = 32'h211ec; force soc.dbg_do = 32'hfec78fa3; #1000;
force soc.dbg_adr = 32'h211f0; force soc.dbg_do = 32'hfee468e3; #1000;
force soc.dbg_adr = 32'h211f4; force soc.dbg_do = 32'h1a050c63; #1000;
force soc.dbg_adr = 32'h211f8; force soc.dbg_do = 32'h3b747463; #1000;
force soc.dbg_adr = 32'h211fc; force soc.dbg_do = 32'h02000693; #1000;
force soc.dbg_adr = 32'h21200; force soc.dbg_do = 32'h03000613; #1000;
force soc.dbg_adr = 32'h21204; force soc.dbg_do = 32'h0cd40a63; #1000;
force soc.dbg_adr = 32'h21208; force soc.dbg_do = 32'h00140413; #1000;
force soc.dbg_adr = 32'h2120c; force soc.dbg_do = 32'h008487b3; #1000;
force soc.dbg_adr = 32'h21210; force soc.dbg_do = 32'hfec78fa3; #1000;
force soc.dbg_adr = 32'h21214; force soc.dbg_do = 32'hff7418e3; #1000;
force soc.dbg_adr = 32'h21218; force soc.dbg_do = 32'hec0598e3; #1000;
force soc.dbg_adr = 32'h2121c; force soc.dbg_do = 32'h000b8713; #1000;
force soc.dbg_adr = 32'h21220; force soc.dbg_do = 32'h00337793; #1000;
force soc.dbg_adr = 32'h21224; force soc.dbg_do = 32'h02000693; #1000;
force soc.dbg_adr = 32'h21228; force soc.dbg_do = 32'heed716e3; #1000;
force soc.dbg_adr = 32'h2122c; force soc.dbg_do = 32'h1c079463; #1000;
force soc.dbg_adr = 32'h21230; force soc.dbg_do = 32'h02000413; #1000;
force soc.dbg_adr = 32'h21234; force soc.dbg_do = 32'hef747ee3; #1000;
force soc.dbg_adr = 32'h21238; force soc.dbg_do = 32'h000b0913; #1000;
force soc.dbg_adr = 32'h2123c; force soc.dbg_do = 32'h41640c33; #1000;
force soc.dbg_adr = 32'h21240; force soc.dbg_do = 32'h00090613; #1000;
force soc.dbg_adr = 32'h21244; force soc.dbg_do = 32'h000a8693; #1000;
force soc.dbg_adr = 32'h21248; force soc.dbg_do = 32'h000a0593; #1000;
force soc.dbg_adr = 32'h2124c; force soc.dbg_do = 32'h02000513; #1000;
force soc.dbg_adr = 32'h21250; force soc.dbg_do = 32'h00190913; #1000;
force soc.dbg_adr = 32'h21254; force soc.dbg_do = 32'h000980e7; #1000;
force soc.dbg_adr = 32'h21258; force soc.dbg_do = 32'h012c07b3; #1000;
force soc.dbg_adr = 32'h2125c; force soc.dbg_do = 32'hff77e2e3; #1000;
force soc.dbg_adr = 32'h21260; force soc.dbg_do = 32'h00140793; #1000;
force soc.dbg_adr = 32'h21264; force soc.dbg_do = 32'h00000c13; #1000;
force soc.dbg_adr = 32'h21268; force soc.dbg_do = 32'h00fbe663; #1000;
force soc.dbg_adr = 32'h2126c; force soc.dbg_do = 32'hfffb8c13; #1000;
force soc.dbg_adr = 32'h21270; force soc.dbg_do = 32'h408c0c33; #1000;
force soc.dbg_adr = 32'h21274; force soc.dbg_do = 32'h001b0793; #1000;
force soc.dbg_adr = 32'h21278; force soc.dbg_do = 32'h00fc0c33; #1000;
force soc.dbg_adr = 32'h2127c; force soc.dbg_do = 32'h0c040c63; #1000;
force soc.dbg_adr = 32'h21280; force soc.dbg_do = 32'h01a12023; #1000;
force soc.dbg_adr = 32'h21284; force soc.dbg_do = 32'heb5ff06f; #1000;
force soc.dbg_adr = 32'h21288; force soc.dbg_do = 32'h08050663; #1000;
force soc.dbg_adr = 32'h2128c; force soc.dbg_do = 32'h16080c63; #1000;
force soc.dbg_adr = 32'h21290; force soc.dbg_do = 32'hfffb8b93; #1000;
force soc.dbg_adr = 32'h21294; force soc.dbg_do = 32'hf4e7e2e3; #1000;
force soc.dbg_adr = 32'h21298; force soc.dbg_do = 32'hf777e2e3; #1000;
force soc.dbg_adr = 32'h2129c; force soc.dbg_do = 32'he40596e3; #1000;
force soc.dbg_adr = 32'h212a0; force soc.dbg_do = 32'h01a12023; #1000;
force soc.dbg_adr = 32'h212a4; force soc.dbg_do = 32'h02000793; #1000;
force soc.dbg_adr = 32'h212a8; force soc.dbg_do = 32'h14f40863; #1000;
force soc.dbg_adr = 32'h212ac; force soc.dbg_do = 32'h0140006f; #1000;
force soc.dbg_adr = 32'h212b0; force soc.dbg_do = 32'h02000793; #1000;
force soc.dbg_adr = 32'h212b4; force soc.dbg_do = 32'he6f40ee3; #1000;
force soc.dbg_adr = 32'h212b8; force soc.dbg_do = 32'h16080c63; #1000;
force soc.dbg_adr = 32'h212bc; force soc.dbg_do = 32'h01a12023; #1000;
force soc.dbg_adr = 32'h212c0; force soc.dbg_do = 32'h008487b3; #1000;
force soc.dbg_adr = 32'h212c4; force soc.dbg_do = 32'h02d00713; #1000;
force soc.dbg_adr = 32'h212c8; force soc.dbg_do = 32'h00e78023; #1000;
force soc.dbg_adr = 32'h212cc; force soc.dbg_do = 32'h00140413; #1000;
force soc.dbg_adr = 32'h212d0; force soc.dbg_do = 32'h000b0c13; #1000;
force soc.dbg_adr = 32'h212d4; force soc.dbg_do = 32'he65ff06f; #1000;
force soc.dbg_adr = 32'h212d8; force soc.dbg_do = 32'h00337793; #1000;
force soc.dbg_adr = 32'h212dc; force soc.dbg_do = 32'hf40588e3; #1000;
force soc.dbg_adr = 32'h212e0; force soc.dbg_do = 32'h40037793; #1000;
force soc.dbg_adr = 32'h212e4; force soc.dbg_do = 32'h08078c63; #1000;
force soc.dbg_adr = 32'h212e8; force soc.dbg_do = 32'h01000713; #1000;
force soc.dbg_adr = 32'h212ec; force soc.dbg_do = 32'h00337793; #1000;
force soc.dbg_adr = 32'h212f0; force soc.dbg_do = 32'h0ce88663; #1000;
force soc.dbg_adr = 32'h212f4; force soc.dbg_do = 32'h00200713; #1000;
force soc.dbg_adr = 32'h212f8; force soc.dbg_do = 32'h06e88263; #1000;
force soc.dbg_adr = 32'h212fc; force soc.dbg_do = 32'h02000713; #1000;
force soc.dbg_adr = 32'h21300; force soc.dbg_do = 32'h16e41e63; #1000;
force soc.dbg_adr = 32'h21304; force soc.dbg_do = 32'he20796e3; #1000;
force soc.dbg_adr = 32'h21308; force soc.dbg_do = 32'he37474e3; #1000;
force soc.dbg_adr = 32'h2130c; force soc.dbg_do = 32'h02000413; #1000;
force soc.dbg_adr = 32'h21310; force soc.dbg_do = 32'hf29ff06f; #1000;
force soc.dbg_adr = 32'h21314; force soc.dbg_do = 32'hece7e2e3; #1000;
force soc.dbg_adr = 32'h21318; force soc.dbg_do = 32'hdc0598e3; #1000;
force soc.dbg_adr = 32'h2131c; force soc.dbg_do = 32'h02000793; #1000;
force soc.dbg_adr = 32'h21320; force soc.dbg_do = 32'hf0f408e3; #1000;
force soc.dbg_adr = 32'h21324; force soc.dbg_do = 32'h00040713; #1000;
force soc.dbg_adr = 32'h21328; force soc.dbg_do = 32'h00337793; #1000;
force soc.dbg_adr = 32'h2132c; force soc.dbg_do = 32'hde0816e3; #1000;
force soc.dbg_adr = 32'h21330; force soc.dbg_do = 32'h00437693; #1000;
force soc.dbg_adr = 32'h21334; force soc.dbg_do = 32'h12068063; #1000;
force soc.dbg_adr = 32'h21338; force soc.dbg_do = 32'h00e486b3; #1000;
force soc.dbg_adr = 32'h2133c; force soc.dbg_do = 32'h02b00613; #1000;
force soc.dbg_adr = 32'h21340; force soc.dbg_do = 32'h00c68023; #1000;
force soc.dbg_adr = 32'h21344; force soc.dbg_do = 32'h00170413; #1000;
force soc.dbg_adr = 32'h21348; force soc.dbg_do = 32'hde0794e3; #1000;
force soc.dbg_adr = 32'h2134c; force soc.dbg_do = 32'hef7466e3; #1000;
force soc.dbg_adr = 32'h21350; force soc.dbg_do = 32'hde1ff06f; #1000;
force soc.dbg_adr = 32'h21354; force soc.dbg_do = 32'h000c0913; #1000;
force soc.dbg_adr = 32'h21358; force soc.dbg_do = 32'he11ff06f; #1000;
force soc.dbg_adr = 32'h2135c; force soc.dbg_do = 32'h02000713; #1000;
force soc.dbg_adr = 32'h21360; force soc.dbg_do = 32'hfae402e3; #1000;
force soc.dbg_adr = 32'h21364; force soc.dbg_do = 32'h00040693; #1000;
force soc.dbg_adr = 32'h21368; force soc.dbg_do = 32'h00140413; #1000;
force soc.dbg_adr = 32'h2136c; force soc.dbg_do = 32'h00d486b3; #1000;
force soc.dbg_adr = 32'h21370; force soc.dbg_do = 32'h06200713; #1000;
force soc.dbg_adr = 32'h21374; force soc.dbg_do = 32'h00e68023; #1000;
force soc.dbg_adr = 32'h21378; force soc.dbg_do = 32'hf85ff06f; #1000;
force soc.dbg_adr = 32'h2137c; force soc.dbg_do = 32'h00870463; #1000;
force soc.dbg_adr = 32'h21380; force soc.dbg_do = 32'hf68b94e3; #1000;
force soc.dbg_adr = 32'h21384; force soc.dbg_do = 32'hfff40693; #1000;
force soc.dbg_adr = 32'h21388; force soc.dbg_do = 32'h01000793; #1000;
force soc.dbg_adr = 32'h2138c; force soc.dbg_do = 32'h10068263; #1000;
force soc.dbg_adr = 32'h21390; force soc.dbg_do = 32'h1ef88663; #1000;
force soc.dbg_adr = 32'h21394; force soc.dbg_do = 32'h00200793; #1000;
force soc.dbg_adr = 32'h21398; force soc.dbg_do = 32'h20f88063; #1000;
force soc.dbg_adr = 32'h2139c; force soc.dbg_do = 32'h00040713; #1000;
force soc.dbg_adr = 32'h213a0; force soc.dbg_do = 32'h00337793; #1000;
force soc.dbg_adr = 32'h213a4; force soc.dbg_do = 32'h00068413; #1000;
force soc.dbg_adr = 32'h213a8; force soc.dbg_do = 32'h0d80006f; #1000;
force soc.dbg_adr = 32'h213ac; force soc.dbg_do = 32'hf2059ae3; #1000;
force soc.dbg_adr = 32'h213b0; force soc.dbg_do = 32'h00040713; #1000;
force soc.dbg_adr = 32'h213b4; force soc.dbg_do = 32'h00337793; #1000;
force soc.dbg_adr = 32'h213b8; force soc.dbg_do = 32'he6dff06f; #1000;
force soc.dbg_adr = 32'h213bc; force soc.dbg_do = 32'h02037713; #1000;
force soc.dbg_adr = 32'h213c0; force soc.dbg_do = 32'h02070063; #1000;
force soc.dbg_adr = 32'h213c4; force soc.dbg_do = 32'h02000713; #1000;
force soc.dbg_adr = 32'h213c8; force soc.dbg_do = 32'h02e40063; #1000;
force soc.dbg_adr = 32'h213cc; force soc.dbg_do = 32'h00848733; #1000;
force soc.dbg_adr = 32'h213d0; force soc.dbg_do = 32'h05800693; #1000;
force soc.dbg_adr = 32'h213d4; force soc.dbg_do = 32'h00d70023; #1000;
force soc.dbg_adr = 32'h213d8; force soc.dbg_do = 32'h00140413; #1000;
force soc.dbg_adr = 32'h213dc; force soc.dbg_do = 32'hf21ff06f; #1000;
force soc.dbg_adr = 32'h213e0; force soc.dbg_do = 32'h02000713; #1000;
force soc.dbg_adr = 32'h213e4; force soc.dbg_do = 32'h10e41a63; #1000;
force soc.dbg_adr = 32'h213e8; force soc.dbg_do = 32'hd40794e3; #1000;
force soc.dbg_adr = 32'h213ec; force soc.dbg_do = 32'he57466e3; #1000;
force soc.dbg_adr = 32'h213f0; force soc.dbg_do = 32'hd41ff06f; #1000;
force soc.dbg_adr = 32'h213f4; force soc.dbg_do = 32'h01a12023; #1000;
force soc.dbg_adr = 32'h213f8; force soc.dbg_do = 32'h000b0c13; #1000;
force soc.dbg_adr = 32'h213fc; force soc.dbg_do = 32'h02000413; #1000;
force soc.dbg_adr = 32'h21400; force soc.dbg_do = 32'hd39ff06f; #1000;
force soc.dbg_adr = 32'h21404; force soc.dbg_do = 32'h00c37793; #1000;
force soc.dbg_adr = 32'h21408; force soc.dbg_do = 32'h00f037b3; #1000;
force soc.dbg_adr = 32'h2140c; force soc.dbg_do = 32'h40fb8bb3; #1000;
force soc.dbg_adr = 32'h21410; force soc.dbg_do = 32'hdce464e3; #1000;
force soc.dbg_adr = 32'h21414; force soc.dbg_do = 32'hdf7464e3; #1000;
force soc.dbg_adr = 32'h21418; force soc.dbg_do = 32'hcc0598e3; #1000;
force soc.dbg_adr = 32'h2141c; force soc.dbg_do = 32'h02000793; #1000;
force soc.dbg_adr = 32'h21420; force soc.dbg_do = 32'hfcf40ae3; #1000;
force soc.dbg_adr = 32'h21424; force soc.dbg_do = 32'h00040713; #1000;
force soc.dbg_adr = 32'h21428; force soc.dbg_do = 32'h00337793; #1000;
force soc.dbg_adr = 32'h2142c; force soc.dbg_do = 32'hf05ff06f; #1000;
force soc.dbg_adr = 32'h21430; force soc.dbg_do = 32'h00437713; #1000;
force soc.dbg_adr = 32'h21434; force soc.dbg_do = 32'h08071263; #1000;
force soc.dbg_adr = 32'h21438; force soc.dbg_do = 32'h00837313; #1000;
force soc.dbg_adr = 32'h2143c; force soc.dbg_do = 32'h10031263; #1000;
force soc.dbg_adr = 32'h21440; force soc.dbg_do = 32'h000b0c13; #1000;
force soc.dbg_adr = 32'h21444; force soc.dbg_do = 32'h000b0913; #1000;
force soc.dbg_adr = 32'h21448; force soc.dbg_do = 32'hd20402e3; #1000;
force soc.dbg_adr = 32'h2144c; force soc.dbg_do = 32'h01a12023; #1000;
force soc.dbg_adr = 32'h21450; force soc.dbg_do = 32'hce9ff06f; #1000;
force soc.dbg_adr = 32'h21454; force soc.dbg_do = 32'h00837313; #1000;
force soc.dbg_adr = 32'h21458; force soc.dbg_do = 32'h06031e63; #1000;
force soc.dbg_adr = 32'h2145c; force soc.dbg_do = 32'h00070413; #1000;
force soc.dbg_adr = 32'h21460; force soc.dbg_do = 32'h10079863; #1000;
force soc.dbg_adr = 32'h21464; force soc.dbg_do = 32'hdd776ae3; #1000;
force soc.dbg_adr = 32'h21468; force soc.dbg_do = 32'h000b0c13; #1000;
force soc.dbg_adr = 32'h2146c; force soc.dbg_do = 32'h000b0913; #1000;
force soc.dbg_adr = 32'h21470; force soc.dbg_do = 32'hd20702e3; #1000;
force soc.dbg_adr = 32'h21474; force soc.dbg_do = 32'h01a12023; #1000;
force soc.dbg_adr = 32'h21478; force soc.dbg_do = 32'hcc1ff06f; #1000;
force soc.dbg_adr = 32'h2147c; force soc.dbg_do = 32'h00140713; #1000;
force soc.dbg_adr = 32'h21480; force soc.dbg_do = 32'h00848433; #1000;
force soc.dbg_adr = 32'h21484; force soc.dbg_do = 32'h03000693; #1000;
force soc.dbg_adr = 32'h21488; force soc.dbg_do = 32'h00d40023; #1000;
force soc.dbg_adr = 32'h2148c; force soc.dbg_do = 32'hd99ff06f; #1000;
force soc.dbg_adr = 32'h21490; force soc.dbg_do = 32'hc6f896e3; #1000;
force soc.dbg_adr = 32'h21494; force soc.dbg_do = 32'h02037793; #1000;
force soc.dbg_adr = 32'h21498; force soc.dbg_do = 32'h0a078063; #1000;
force soc.dbg_adr = 32'h2149c; force soc.dbg_do = 32'h05800713; #1000;
force soc.dbg_adr = 32'h214a0; force soc.dbg_do = 32'h03000793; #1000;
force soc.dbg_adr = 32'h214a4; force soc.dbg_do = 32'h00e48023; #1000;
force soc.dbg_adr = 32'h214a8; force soc.dbg_do = 32'h00f480a3; #1000;
force soc.dbg_adr = 32'h214ac; force soc.dbg_do = 32'h00200713; #1000;
force soc.dbg_adr = 32'h214b0; force soc.dbg_do = 32'h00337793; #1000;
force soc.dbg_adr = 32'h214b4; force soc.dbg_do = 32'hc61ff06f; #1000;
force soc.dbg_adr = 32'h214b8; force soc.dbg_do = 32'h008487b3; #1000;
force soc.dbg_adr = 32'h214bc; force soc.dbg_do = 32'h01a12023; #1000;
force soc.dbg_adr = 32'h214c0; force soc.dbg_do = 32'h02b00713; #1000;
force soc.dbg_adr = 32'h214c4; force soc.dbg_do = 32'h00e78023; #1000;
force soc.dbg_adr = 32'h214c8; force soc.dbg_do = 32'h00140413; #1000;
force soc.dbg_adr = 32'h214cc; force soc.dbg_do = 32'h000b0c13; #1000;
force soc.dbg_adr = 32'h214d0; force soc.dbg_do = 32'hc69ff06f; #1000;
force soc.dbg_adr = 32'h214d4; force soc.dbg_do = 32'h00e486b3; #1000;
force soc.dbg_adr = 32'h214d8; force soc.dbg_do = 32'h02000613; #1000;
force soc.dbg_adr = 32'h214dc; force soc.dbg_do = 32'h00c68023; #1000;
force soc.dbg_adr = 32'h214e0; force soc.dbg_do = 32'h00170413; #1000;
force soc.dbg_adr = 32'h214e4; force soc.dbg_do = 32'hf00784e3; #1000;
force soc.dbg_adr = 32'h214e8; force soc.dbg_do = 32'hc49ff06f; #1000;
force soc.dbg_adr = 32'h214ec; force soc.dbg_do = 32'h01a12023; #1000;
force soc.dbg_adr = 32'h214f0; force soc.dbg_do = 32'h000b0c13; #1000;
force soc.dbg_adr = 32'h214f4; force soc.dbg_do = 32'hc45ff06f; #1000;
force soc.dbg_adr = 32'h214f8; force soc.dbg_do = 32'h00848733; #1000;
force soc.dbg_adr = 32'h214fc; force soc.dbg_do = 32'h07800693; #1000;
force soc.dbg_adr = 32'h21500; force soc.dbg_do = 32'h00d70023; #1000;
force soc.dbg_adr = 32'h21504; force soc.dbg_do = 32'h00140413; #1000;
force soc.dbg_adr = 32'h21508; force soc.dbg_do = 32'hdf5ff06f; #1000;
force soc.dbg_adr = 32'h2150c; force soc.dbg_do = 32'h02037793; #1000;
force soc.dbg_adr = 32'h21510; force soc.dbg_do = 32'h02078463; #1000;
force soc.dbg_adr = 32'h21514; force soc.dbg_do = 32'h05800793; #1000;
force soc.dbg_adr = 32'h21518; force soc.dbg_do = 32'h03000713; #1000;
force soc.dbg_adr = 32'h2151c; force soc.dbg_do = 32'h00f48023; #1000;
force soc.dbg_adr = 32'h21520; force soc.dbg_do = 32'h00e480a3; #1000;
force soc.dbg_adr = 32'h21524; force soc.dbg_do = 32'h00337793; #1000;
force soc.dbg_adr = 32'h21528; force soc.dbg_do = 32'h00200713; #1000;
force soc.dbg_adr = 32'h2152c; force soc.dbg_do = 32'hbe9ff06f; #1000;
force soc.dbg_adr = 32'h21530; force soc.dbg_do = 32'h06200793; #1000;
force soc.dbg_adr = 32'h21534; force soc.dbg_do = 32'hfe5ff06f; #1000;
force soc.dbg_adr = 32'h21538; force soc.dbg_do = 32'h07800793; #1000;
force soc.dbg_adr = 32'h2153c; force soc.dbg_do = 32'hfddff06f; #1000;
force soc.dbg_adr = 32'h21540; force soc.dbg_do = 32'h00848733; #1000;
force soc.dbg_adr = 32'h21544; force soc.dbg_do = 32'h01a12023; #1000;
force soc.dbg_adr = 32'h21548; force soc.dbg_do = 32'h00f70023; #1000;
force soc.dbg_adr = 32'h2154c; force soc.dbg_do = 32'h00140413; #1000;
force soc.dbg_adr = 32'h21550; force soc.dbg_do = 32'h000b0c13; #1000;
force soc.dbg_adr = 32'h21554; force soc.dbg_do = 32'hbe5ff06f; #1000;
force soc.dbg_adr = 32'h21558; force soc.dbg_do = 32'h04058663; #1000;
force soc.dbg_adr = 32'h2155c; force soc.dbg_do = 32'h40037793; #1000;
force soc.dbg_adr = 32'h21560; force soc.dbg_do = 32'hd80794e3; #1000;
force soc.dbg_adr = 32'h21564; force soc.dbg_do = 32'hb80408e3; #1000;
force soc.dbg_adr = 32'h21568; force soc.dbg_do = 32'hd8e410e3; #1000;
force soc.dbg_adr = 32'h2156c; force soc.dbg_do = 32'he19ff06f; #1000;
force soc.dbg_adr = 32'h21570; force soc.dbg_do = 32'h000b0c13; #1000;
force soc.dbg_adr = 32'h21574; force soc.dbg_do = 32'hd00416e3; #1000;
force soc.dbg_adr = 32'h21578; force soc.dbg_do = 32'hdddff06f; #1000;
force soc.dbg_adr = 32'h2157c; force soc.dbg_do = 32'hffe40793; #1000;
force soc.dbg_adr = 32'h21580; force soc.dbg_do = 32'h02037713; #1000;
force soc.dbg_adr = 32'h21584; force soc.dbg_do = 32'h00f487b3; #1000;
force soc.dbg_adr = 32'h21588; force soc.dbg_do = 32'h02070463; #1000;
force soc.dbg_adr = 32'h2158c; force soc.dbg_do = 32'h05800713; #1000;
force soc.dbg_adr = 32'h21590; force soc.dbg_do = 32'h00e78023; #1000;
force soc.dbg_adr = 32'h21594; force soc.dbg_do = 32'he09ff06f; #1000;
force soc.dbg_adr = 32'h21598; force soc.dbg_do = 32'h00337793; #1000;
force soc.dbg_adr = 32'h2159c; force soc.dbg_do = 32'hdd1ff06f; #1000;
force soc.dbg_adr = 32'h215a0; force soc.dbg_do = 32'hd40590e3; #1000;
force soc.dbg_adr = 32'h215a4; force soc.dbg_do = 32'h02000793; #1000;
force soc.dbg_adr = 32'h215a8; force soc.dbg_do = 32'hb8f404e3; #1000;
force soc.dbg_adr = 32'h215ac; force soc.dbg_do = 32'hd79ff06f; #1000;
force soc.dbg_adr = 32'h215b0; force soc.dbg_do = 32'h07800713; #1000;
force soc.dbg_adr = 32'h215b4; force soc.dbg_do = 32'h00e78023; #1000;
force soc.dbg_adr = 32'h215b8; force soc.dbg_do = 32'hde5ff06f; #1000;
force soc.dbg_adr = 32'h215bc; force soc.dbg_do = 32'h00051463; #1000;
force soc.dbg_adr = 32'h215c0; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h215c4; force soc.dbg_do = 32'ha79fe06f; #1000;
force soc.dbg_adr = 32'h215c8; force soc.dbg_do = 32'h00050863; #1000;
force soc.dbg_adr = 32'h215cc; force soc.dbg_do = 32'h0005a783; #1000;
force soc.dbg_adr = 32'h215d0; force soc.dbg_do = 32'h0045a583; #1000;
force soc.dbg_adr = 32'h215d4; force soc.dbg_do = 32'h00078067; #1000;
force soc.dbg_adr = 32'h215d8; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h215dc; force soc.dbg_do = 32'hf6010113; #1000;
force soc.dbg_adr = 32'h215e0; force soc.dbg_do = 32'h08912a23; #1000;
force soc.dbg_adr = 32'h215e4; force soc.dbg_do = 32'h09312623; #1000;
force soc.dbg_adr = 32'h215e8; force soc.dbg_do = 32'h07812c23; #1000;
force soc.dbg_adr = 32'h215ec; force soc.dbg_do = 32'h07b12623; #1000;
force soc.dbg_adr = 32'h215f0; force soc.dbg_do = 32'h08112e23; #1000;
force soc.dbg_adr = 32'h215f4; force soc.dbg_do = 32'h08812c23; #1000;
force soc.dbg_adr = 32'h215f8; force soc.dbg_do = 32'h07712e23; #1000;
force soc.dbg_adr = 32'h215fc; force soc.dbg_do = 32'h00b12c23; #1000;
force soc.dbg_adr = 32'h21600; force soc.dbg_do = 32'h00060493; #1000;
force soc.dbg_adr = 32'h21604; force soc.dbg_do = 32'h00068c13; #1000;
force soc.dbg_adr = 32'h21608; force soc.dbg_do = 32'h00070d93; #1000;
force soc.dbg_adr = 32'h2160c; force soc.dbg_do = 32'h00050993; #1000;
force soc.dbg_adr = 32'h21610; force soc.dbg_do = 32'h64058663; #1000;
force soc.dbg_adr = 32'h21614; force soc.dbg_do = 32'h000c4503; #1000;
force soc.dbg_adr = 32'h21618; force soc.dbg_do = 32'h00000b93; #1000;
force soc.dbg_adr = 32'h2161c; force soc.dbg_do = 32'h64050a63; #1000;
force soc.dbg_adr = 32'h21620; force soc.dbg_do = 32'h000c0793; #1000;
force soc.dbg_adr = 32'h21624; force soc.dbg_do = 32'h09412423; #1000;
force soc.dbg_adr = 32'h21628; force soc.dbg_do = 32'h09512223; #1000;
force soc.dbg_adr = 32'h2162c; force soc.dbg_do = 32'h09612023; #1000;
force soc.dbg_adr = 32'h21630; force soc.dbg_do = 32'h000b8c13; #1000;
force soc.dbg_adr = 32'h21634; force soc.dbg_do = 32'h09212823; #1000;
force soc.dbg_adr = 32'h21638; force soc.dbg_do = 32'h07912a23; #1000;
force soc.dbg_adr = 32'h2163c; force soc.dbg_do = 32'h02500b13; #1000;
force soc.dbg_adr = 32'h21640; force soc.dbg_do = 32'h01000413; #1000;
force soc.dbg_adr = 32'h21644; force soc.dbg_do = 32'h00024a37; #1000;
force soc.dbg_adr = 32'h21648; force soc.dbg_do = 32'h00900a93; #1000;
force soc.dbg_adr = 32'h2164c; force soc.dbg_do = 32'h00078b93; #1000;
force soc.dbg_adr = 32'h21650; force soc.dbg_do = 32'h0200006f; #1000;
force soc.dbg_adr = 32'h21654; force soc.dbg_do = 32'h01812583; #1000;
force soc.dbg_adr = 32'h21658; force soc.dbg_do = 32'h000c0613; #1000;
force soc.dbg_adr = 32'h2165c; force soc.dbg_do = 32'h00048693; #1000;
force soc.dbg_adr = 32'h21660; force soc.dbg_do = 32'h001c0c13; #1000;
force soc.dbg_adr = 32'h21664; force soc.dbg_do = 32'h000980e7; #1000;
force soc.dbg_adr = 32'h21668; force soc.dbg_do = 32'h000bc503; #1000;
force soc.dbg_adr = 32'h2166c; force soc.dbg_do = 32'h22050a63; #1000;
force soc.dbg_adr = 32'h21670; force soc.dbg_do = 32'h001b8b93; #1000;
force soc.dbg_adr = 32'h21674; force soc.dbg_do = 32'hff6510e3; #1000;
force soc.dbg_adr = 32'h21678; force soc.dbg_do = 32'h00000693; #1000;
force soc.dbg_adr = 32'h2167c; force soc.dbg_do = 32'h000bc503; #1000;
force soc.dbg_adr = 32'h21680; force soc.dbg_do = 32'h001b8713; #1000;
force soc.dbg_adr = 32'h21684; force soc.dbg_do = 32'hfe050793; #1000;
force soc.dbg_adr = 32'h21688; force soc.dbg_do = 32'h0ff7f793; #1000;
force soc.dbg_adr = 32'h2168c; force soc.dbg_do = 32'h00f46c63; #1000;
force soc.dbg_adr = 32'h21690; force soc.dbg_do = 32'h00279793; #1000;
force soc.dbg_adr = 32'h21694; force soc.dbg_do = 32'h13ca0613; #1000;
force soc.dbg_adr = 32'h21698; force soc.dbg_do = 32'h00c787b3; #1000;
force soc.dbg_adr = 32'h2169c; force soc.dbg_do = 32'h0007a783; #1000;
force soc.dbg_adr = 32'h216a0; force soc.dbg_do = 32'h00078067; #1000;
force soc.dbg_adr = 32'h216a4; force soc.dbg_do = 32'hfd050793; #1000;
force soc.dbg_adr = 32'h216a8; force soc.dbg_do = 32'h0ff7f793; #1000;
force soc.dbg_adr = 32'h216ac; force soc.dbg_do = 32'h24fafa63; #1000;
force soc.dbg_adr = 32'h216b0; force soc.dbg_do = 32'h02a00793; #1000;
force soc.dbg_adr = 32'h216b4; force soc.dbg_do = 32'h00000e13; #1000;
force soc.dbg_adr = 32'h216b8; force soc.dbg_do = 32'h2cf50263; #1000;
force soc.dbg_adr = 32'h216bc; force soc.dbg_do = 32'h02e00793; #1000;
force soc.dbg_adr = 32'h216c0; force soc.dbg_do = 32'h00000e93; #1000;
force soc.dbg_adr = 32'h216c4; force soc.dbg_do = 32'h28f50463; #1000;
force soc.dbg_adr = 32'h216c8; force soc.dbg_do = 32'hf9850793; #1000;
force soc.dbg_adr = 32'h216cc; force soc.dbg_do = 32'h0ff7f793; #1000;
force soc.dbg_adr = 32'h216d0; force soc.dbg_do = 32'h01200613; #1000;
force soc.dbg_adr = 32'h216d4; force soc.dbg_do = 32'h06f66263; #1000;
force soc.dbg_adr = 32'h216d8; force soc.dbg_do = 32'h00024637; #1000;
force soc.dbg_adr = 32'h216dc; force soc.dbg_do = 32'h00279793; #1000;
force soc.dbg_adr = 32'h216e0; force soc.dbg_do = 32'h18060613; #1000;
force soc.dbg_adr = 32'h216e4; force soc.dbg_do = 32'h00c787b3; #1000;
force soc.dbg_adr = 32'h216e8; force soc.dbg_do = 32'h0007a783; #1000;
force soc.dbg_adr = 32'h216ec; force soc.dbg_do = 32'h00078067; #1000;
force soc.dbg_adr = 32'h216f0; force soc.dbg_do = 32'h0016e693; #1000;
force soc.dbg_adr = 32'h216f4; force soc.dbg_do = 32'h00070b93; #1000;
force soc.dbg_adr = 32'h216f8; force soc.dbg_do = 32'hf85ff06f; #1000;
force soc.dbg_adr = 32'h216fc; force soc.dbg_do = 32'h0026e693; #1000;
force soc.dbg_adr = 32'h21700; force soc.dbg_do = 32'h00070b93; #1000;
force soc.dbg_adr = 32'h21704; force soc.dbg_do = 32'hf79ff06f; #1000;
force soc.dbg_adr = 32'h21708; force soc.dbg_do = 32'h0046e693; #1000;
force soc.dbg_adr = 32'h2170c; force soc.dbg_do = 32'h00070b93; #1000;
force soc.dbg_adr = 32'h21710; force soc.dbg_do = 32'hf6dff06f; #1000;
force soc.dbg_adr = 32'h21714; force soc.dbg_do = 32'h0106e693; #1000;
force soc.dbg_adr = 32'h21718; force soc.dbg_do = 32'h00070b93; #1000;
force soc.dbg_adr = 32'h2171c; force soc.dbg_do = 32'hf61ff06f; #1000;
force soc.dbg_adr = 32'h21720; force soc.dbg_do = 32'h0086e693; #1000;
force soc.dbg_adr = 32'h21724; force soc.dbg_do = 32'h00070b93; #1000;
force soc.dbg_adr = 32'h21728; force soc.dbg_do = 32'hf55ff06f; #1000;
force soc.dbg_adr = 32'h2172c; force soc.dbg_do = 32'h001bc503; #1000;
force soc.dbg_adr = 32'h21730; force soc.dbg_do = 32'h1006e693; #1000;
force soc.dbg_adr = 32'h21734; force soc.dbg_do = 32'h00170713; #1000;
force soc.dbg_adr = 32'h21738; force soc.dbg_do = 32'h07800613; #1000;
force soc.dbg_adr = 32'h2173c; force soc.dbg_do = 32'h00070b93; #1000;
force soc.dbg_adr = 32'h21740; force soc.dbg_do = 32'hf0a66ae3; #1000;
force soc.dbg_adr = 32'h21744; force soc.dbg_do = 32'h06300793; #1000;
force soc.dbg_adr = 32'h21748; force soc.dbg_do = 32'h0aa7e063; #1000;
force soc.dbg_adr = 32'h2174c; force soc.dbg_do = 32'h06200713; #1000;
force soc.dbg_adr = 32'h21750; force soc.dbg_do = 32'h72e50863; #1000;
force soc.dbg_adr = 32'h21754; force soc.dbg_do = 32'h36f50a63; #1000;
force soc.dbg_adr = 32'h21758; force soc.dbg_do = 32'h02500793; #1000;
force soc.dbg_adr = 32'h2175c; force soc.dbg_do = 32'heef50ce3; #1000;
force soc.dbg_adr = 32'h21760; force soc.dbg_do = 32'h05800793; #1000;
force soc.dbg_adr = 32'h21764; force soc.dbg_do = 32'heef518e3; #1000;
force soc.dbg_adr = 32'h21768; force soc.dbg_do = 32'h01000613; #1000;
force soc.dbg_adr = 32'h2176c; force soc.dbg_do = 32'h07a12823; #1000;
force soc.dbg_adr = 32'h21770; force soc.dbg_do = 32'h0206e693; #1000;
force soc.dbg_adr = 32'h21774; force soc.dbg_do = 32'h00060893; #1000;
force soc.dbg_adr = 32'h21778; force soc.dbg_do = 32'h00000f13; #1000;
force soc.dbg_adr = 32'h2177c; force soc.dbg_do = 32'h4006f593; #1000;
force soc.dbg_adr = 32'h21780; force soc.dbg_do = 32'hff36f813; #1000;
force soc.dbg_adr = 32'h21784; force soc.dbg_do = 32'h00058463; #1000;
force soc.dbg_adr = 32'h21788; force soc.dbg_do = 32'hff26f813; #1000;
force soc.dbg_adr = 32'h2178c; force soc.dbg_do = 32'h20087c93; #1000;
force soc.dbg_adr = 32'h21790; force soc.dbg_do = 32'h700c9263; #1000;
force soc.dbg_adr = 32'h21794; force soc.dbg_do = 32'h004d8793; #1000;
force soc.dbg_adr = 32'h21798; force soc.dbg_do = 32'h10087d13; #1000;
force soc.dbg_adr = 32'h2179c; force soc.dbg_do = 32'h00f12e23; #1000;
force soc.dbg_adr = 32'h217a0; force soc.dbg_do = 32'h400d1ce3; #1000;
force soc.dbg_adr = 32'h217a4; force soc.dbg_do = 32'h04087793; #1000;
force soc.dbg_adr = 32'h217a8; force soc.dbg_do = 32'h060794e3; #1000;
force soc.dbg_adr = 32'h217ac; force soc.dbg_do = 32'h08087793; #1000;
force soc.dbg_adr = 32'h217b0; force soc.dbg_do = 32'h520782e3; #1000;
force soc.dbg_adr = 32'h217b4; force soc.dbg_do = 32'h000ddc83; #1000;
force soc.dbg_adr = 32'h217b8; force soc.dbg_do = 32'h220c98e3; #1000;
force soc.dbg_adr = 32'h217bc; force soc.dbg_do = 32'hfef87813; #1000;
force soc.dbg_adr = 32'h217c0; force soc.dbg_do = 32'h220584e3; #1000;
force soc.dbg_adr = 32'h217c4; force soc.dbg_do = 32'h00000d13; #1000;
force soc.dbg_adr = 32'h217c8; force soc.dbg_do = 32'h04010713; #1000;
force soc.dbg_adr = 32'h217cc; force soc.dbg_do = 32'h01012423; #1000;
force soc.dbg_adr = 32'h217d0; force soc.dbg_do = 32'h01c12223; #1000;
force soc.dbg_adr = 32'h217d4; force soc.dbg_do = 32'h01d12023; #1000;
force soc.dbg_adr = 32'h217d8; force soc.dbg_do = 32'h000d0793; #1000;
force soc.dbg_adr = 32'h217dc; force soc.dbg_do = 32'h000c0613; #1000;
force soc.dbg_adr = 32'h217e0; force soc.dbg_do = 32'h00000813; #1000;
force soc.dbg_adr = 32'h217e4; force soc.dbg_do = 32'h4580006f; #1000;
force soc.dbg_adr = 32'h217e8; force soc.dbg_do = 32'hf9c50713; #1000;
force soc.dbg_adr = 32'h217ec; force soc.dbg_do = 32'h00100c93; #1000;
force soc.dbg_adr = 32'h217f0; force soc.dbg_do = 32'h001217b7; #1000;
force soc.dbg_adr = 32'h217f4; force soc.dbg_do = 32'h00ec9cb3; #1000;
force soc.dbg_adr = 32'h217f8; force soc.dbg_do = 32'h82178793; #1000;
force soc.dbg_adr = 32'h217fc; force soc.dbg_do = 32'h00fcfcb3; #1000;
force soc.dbg_adr = 32'h21800; force soc.dbg_do = 32'h320c9863; #1000;
force soc.dbg_adr = 32'h21804; force soc.dbg_do = 32'h07300793; #1000;
force soc.dbg_adr = 32'h21808; force soc.dbg_do = 32'h1ef50663; #1000;
force soc.dbg_adr = 32'h2180c; force soc.dbg_do = 32'h07000793; #1000;
force soc.dbg_adr = 32'h21810; force soc.dbg_do = 32'he4f512e3; #1000;
force soc.dbg_adr = 32'h21814; force soc.dbg_do = 32'h000da783; #1000;
force soc.dbg_adr = 32'h21818; force soc.dbg_do = 32'h0216e613; #1000;
force soc.dbg_adr = 32'h2181c; force soc.dbg_do = 32'h004d8d93; #1000;
force soc.dbg_adr = 32'h21820; force soc.dbg_do = 32'h4a078c63; #1000;
force soc.dbg_adr = 32'h21824; force soc.dbg_do = 32'h04010713; #1000;
force soc.dbg_adr = 32'h21828; force soc.dbg_do = 32'h00900813; #1000;
force soc.dbg_adr = 32'h2182c; force soc.dbg_do = 32'h00f00513; #1000;
force soc.dbg_adr = 32'h21830; force soc.dbg_do = 32'h02000893; #1000;
force soc.dbg_adr = 32'h21834; force soc.dbg_do = 32'h00c0006f; #1000;
force soc.dbg_adr = 32'h21838; force soc.dbg_do = 32'h031c8663; #1000;
force soc.dbg_adr = 32'h2183c; force soc.dbg_do = 32'h00068793; #1000;
force soc.dbg_adr = 32'h21840; force soc.dbg_do = 32'h00f7f313; #1000;
force soc.dbg_adr = 32'h21844; force soc.dbg_do = 32'h03730593; #1000;
force soc.dbg_adr = 32'h21848; force soc.dbg_do = 32'h00686463; #1000;
force soc.dbg_adr = 32'h2184c; force soc.dbg_do = 32'h03030593; #1000;
force soc.dbg_adr = 32'h21850; force soc.dbg_do = 32'h001c8c93; #1000;
force soc.dbg_adr = 32'h21854; force soc.dbg_do = 32'h019706b3; #1000;
force soc.dbg_adr = 32'h21858; force soc.dbg_do = 32'hfeb68fa3; #1000;
force soc.dbg_adr = 32'h2185c; force soc.dbg_do = 32'h0047d693; #1000;
force soc.dbg_adr = 32'h21860; force soc.dbg_do = 32'hfcf56ce3; #1000;
force soc.dbg_adr = 32'h21864; force soc.dbg_do = 32'h01812583; #1000;
force soc.dbg_adr = 32'h21868; force soc.dbg_do = 32'h00800693; #1000;
force soc.dbg_adr = 32'h2186c; force soc.dbg_do = 32'h00c12423; #1000;
force soc.dbg_adr = 32'h21870; force soc.dbg_do = 32'h00d12223; #1000;
force soc.dbg_adr = 32'h21874; force soc.dbg_do = 32'h000c0613; #1000;
force soc.dbg_adr = 32'h21878; force soc.dbg_do = 32'h01d12023; #1000;
force soc.dbg_adr = 32'h2187c; force soc.dbg_do = 32'h000c8793; #1000;
force soc.dbg_adr = 32'h21880; force soc.dbg_do = 32'h01000893; #1000;
force soc.dbg_adr = 32'h21884; force soc.dbg_do = 32'h00000813; #1000;
force soc.dbg_adr = 32'h21888; force soc.dbg_do = 32'h00048693; #1000;
force soc.dbg_adr = 32'h2188c; force soc.dbg_do = 32'h00098513; #1000;
force soc.dbg_adr = 32'h21890; force soc.dbg_do = 32'hff4ff0ef; #1000;
force soc.dbg_adr = 32'h21894; force soc.dbg_do = 32'h00050c13; #1000;
force soc.dbg_adr = 32'h21898; force soc.dbg_do = 32'h000bc503; #1000;
force soc.dbg_adr = 32'h2189c; force soc.dbg_do = 32'hdc051ae3; #1000;
force soc.dbg_adr = 32'h218a0; force soc.dbg_do = 32'h000c0b93; #1000;
force soc.dbg_adr = 32'h218a4; force soc.dbg_do = 32'h09012903; #1000;
force soc.dbg_adr = 32'h218a8; force soc.dbg_do = 32'h08812a03; #1000;
force soc.dbg_adr = 32'h218ac; force soc.dbg_do = 32'h08412a83; #1000;
force soc.dbg_adr = 32'h218b0; force soc.dbg_do = 32'h08012b03; #1000;
force soc.dbg_adr = 32'h218b4; force soc.dbg_do = 32'h07412c83; #1000;
force soc.dbg_adr = 32'h218b8; force soc.dbg_do = 32'h000c0413; #1000;
force soc.dbg_adr = 32'h218bc; force soc.dbg_do = 32'h009be463; #1000;
force soc.dbg_adr = 32'h218c0; force soc.dbg_do = 32'hfff48b93; #1000;
force soc.dbg_adr = 32'h218c4; force soc.dbg_do = 32'h01812583; #1000;
force soc.dbg_adr = 32'h218c8; force soc.dbg_do = 32'h00048693; #1000;
force soc.dbg_adr = 32'h218cc; force soc.dbg_do = 32'h000b8613; #1000;
force soc.dbg_adr = 32'h218d0; force soc.dbg_do = 32'h00000513; #1000;
force soc.dbg_adr = 32'h218d4; force soc.dbg_do = 32'h000980e7; #1000;
force soc.dbg_adr = 32'h218d8; force soc.dbg_do = 32'h09c12083; #1000;
force soc.dbg_adr = 32'h218dc; force soc.dbg_do = 32'h00040513; #1000;
force soc.dbg_adr = 32'h218e0; force soc.dbg_do = 32'h09812403; #1000;
force soc.dbg_adr = 32'h218e4; force soc.dbg_do = 32'h09412483; #1000;
force soc.dbg_adr = 32'h218e8; force soc.dbg_do = 32'h08c12983; #1000;
force soc.dbg_adr = 32'h218ec; force soc.dbg_do = 32'h07c12b83; #1000;
force soc.dbg_adr = 32'h218f0; force soc.dbg_do = 32'h07812c03; #1000;
force soc.dbg_adr = 32'h218f4; force soc.dbg_do = 32'h06c12d83; #1000;
force soc.dbg_adr = 32'h218f8; force soc.dbg_do = 32'h0a010113; #1000;
force soc.dbg_adr = 32'h218fc; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h21900; force soc.dbg_do = 32'h00000e13; #1000;
force soc.dbg_adr = 32'h21904; force soc.dbg_do = 32'h000e0613; #1000;
force soc.dbg_adr = 32'h21908; force soc.dbg_do = 32'h0080006f; #1000;
force soc.dbg_adr = 32'h2190c; force soc.dbg_do = 32'h00170713; #1000;
force soc.dbg_adr = 32'h21910; force soc.dbg_do = 32'h00261e13; #1000;
force soc.dbg_adr = 32'h21914; force soc.dbg_do = 32'h00ce0e33; #1000;
force soc.dbg_adr = 32'h21918; force soc.dbg_do = 32'h001e1e13; #1000;
force soc.dbg_adr = 32'h2191c; force soc.dbg_do = 32'h00ae0e33; #1000;
force soc.dbg_adr = 32'h21920; force soc.dbg_do = 32'h00074503; #1000;
force soc.dbg_adr = 32'h21924; force soc.dbg_do = 32'hfd0e0613; #1000;
force soc.dbg_adr = 32'h21928; force soc.dbg_do = 32'h00070b93; #1000;
force soc.dbg_adr = 32'h2192c; force soc.dbg_do = 32'hfd050793; #1000;
force soc.dbg_adr = 32'h21930; force soc.dbg_do = 32'h0ff7f793; #1000;
force soc.dbg_adr = 32'h21934; force soc.dbg_do = 32'hfcfafce3; #1000;
force soc.dbg_adr = 32'h21938; force soc.dbg_do = 32'h02e00793; #1000;
force soc.dbg_adr = 32'h2193c; force soc.dbg_do = 32'h00060e13; #1000;
force soc.dbg_adr = 32'h21940; force soc.dbg_do = 32'h00170713; #1000;
force soc.dbg_adr = 32'h21944; force soc.dbg_do = 32'h00000e93; #1000;
force soc.dbg_adr = 32'h21948; force soc.dbg_do = 32'hd8f510e3; #1000;
force soc.dbg_adr = 32'h2194c; force soc.dbg_do = 32'h001bc503; #1000;
force soc.dbg_adr = 32'h21950; force soc.dbg_do = 32'h00900793; #1000;
force soc.dbg_adr = 32'h21954; force soc.dbg_do = 32'h4006e693; #1000;
force soc.dbg_adr = 32'h21958; force soc.dbg_do = 32'hfd050593; #1000;
force soc.dbg_adr = 32'h2195c; force soc.dbg_do = 32'h0ff5f593; #1000;
force soc.dbg_adr = 32'h21960; force soc.dbg_do = 32'h00070613; #1000;
force soc.dbg_adr = 32'h21964; force soc.dbg_do = 32'h30b7fc63; #1000;
force soc.dbg_adr = 32'h21968; force soc.dbg_do = 32'h02a00793; #1000;
force soc.dbg_adr = 32'h2196c; force soc.dbg_do = 32'h34f50463; #1000;
force soc.dbg_adr = 32'h21970; force soc.dbg_do = 32'h00070b93; #1000;
force soc.dbg_adr = 32'h21974; force soc.dbg_do = 32'h00170713; #1000;
force soc.dbg_adr = 32'h21978; force soc.dbg_do = 32'hd51ff06f; #1000;
force soc.dbg_adr = 32'h2197c; force soc.dbg_do = 32'h000dae03; #1000;
force soc.dbg_adr = 32'h21980; force soc.dbg_do = 32'h004d8d93; #1000;
force soc.dbg_adr = 32'h21984; force soc.dbg_do = 32'h000e4a63; #1000;
force soc.dbg_adr = 32'h21988; force soc.dbg_do = 32'h001bc503; #1000;
force soc.dbg_adr = 32'h2198c; force soc.dbg_do = 32'h00070b93; #1000;
force soc.dbg_adr = 32'h21990; force soc.dbg_do = 32'h00170713; #1000;
force soc.dbg_adr = 32'h21994; force soc.dbg_do = 32'hd29ff06f; #1000;
force soc.dbg_adr = 32'h21998; force soc.dbg_do = 32'h001bc503; #1000;
force soc.dbg_adr = 32'h2199c; force soc.dbg_do = 32'h0026e693; #1000;
force soc.dbg_adr = 32'h219a0; force soc.dbg_do = 32'h00070b93; #1000;
force soc.dbg_adr = 32'h219a4; force soc.dbg_do = 32'h41c00e33; #1000;
force soc.dbg_adr = 32'h219a8; force soc.dbg_do = 32'h00170713; #1000;
force soc.dbg_adr = 32'h219ac; force soc.dbg_do = 32'hd11ff06f; #1000;
force soc.dbg_adr = 32'h219b0; force soc.dbg_do = 32'h001bc503; #1000;
force soc.dbg_adr = 32'h219b4; force soc.dbg_do = 32'h06c00793; #1000;
force soc.dbg_adr = 32'h219b8; force soc.dbg_do = 32'hd6f51ce3; #1000;
force soc.dbg_adr = 32'h219bc; force soc.dbg_do = 32'h002bc503; #1000;
force soc.dbg_adr = 32'h219c0; force soc.dbg_do = 32'h3006e693; #1000;
force soc.dbg_adr = 32'h219c4; force soc.dbg_do = 32'h003b8713; #1000;
force soc.dbg_adr = 32'h219c8; force soc.dbg_do = 32'hd71ff06f; #1000;
force soc.dbg_adr = 32'h219cc; force soc.dbg_do = 32'h001bc503; #1000;
force soc.dbg_adr = 32'h219d0; force soc.dbg_do = 32'h2006e693; #1000;
force soc.dbg_adr = 32'h219d4; force soc.dbg_do = 32'h00170713; #1000;
force soc.dbg_adr = 32'h219d8; force soc.dbg_do = 32'hd61ff06f; #1000;
force soc.dbg_adr = 32'h219dc; force soc.dbg_do = 32'h001bc503; #1000;
force soc.dbg_adr = 32'h219e0; force soc.dbg_do = 32'h06800793; #1000;
force soc.dbg_adr = 32'h219e4; force soc.dbg_do = 32'h3af50063; #1000;
force soc.dbg_adr = 32'h219e8; force soc.dbg_do = 32'h0806e693; #1000;
force soc.dbg_adr = 32'h219ec; force soc.dbg_do = 32'h00170713; #1000;
force soc.dbg_adr = 32'h219f0; force soc.dbg_do = 32'hd49ff06f; #1000;
force soc.dbg_adr = 32'h219f4; force soc.dbg_do = 32'h07a12823; #1000;
force soc.dbg_adr = 32'h219f8; force soc.dbg_do = 32'h004d8913; #1000;
force soc.dbg_adr = 32'h219fc; force soc.dbg_do = 32'hfff00613; #1000;
force soc.dbg_adr = 32'h21a00; force soc.dbg_do = 32'h000dad83; #1000;
force soc.dbg_adr = 32'h21a04; force soc.dbg_do = 32'h000e8463; #1000;
force soc.dbg_adr = 32'h21a08; force soc.dbg_do = 32'h000e8613; #1000;
force soc.dbg_adr = 32'h21a0c; force soc.dbg_do = 32'h000dc503; #1000;
force soc.dbg_adr = 32'h21a10; force soc.dbg_do = 32'h00cd8633; #1000;
force soc.dbg_adr = 32'h21a14; force soc.dbg_do = 32'h000d8793; #1000;
force soc.dbg_adr = 32'h21a18; force soc.dbg_do = 32'h40050a63; #1000;
force soc.dbg_adr = 32'h21a1c; force soc.dbg_do = 32'h2ef60663; #1000;
force soc.dbg_adr = 32'h21a20; force soc.dbg_do = 32'h0017c703; #1000;
force soc.dbg_adr = 32'h21a24; force soc.dbg_do = 32'h00178793; #1000;
force soc.dbg_adr = 32'h21a28; force soc.dbg_do = 32'hfe071ae3; #1000;
force soc.dbg_adr = 32'h21a2c; force soc.dbg_do = 32'h4006f713; #1000;
force soc.dbg_adr = 32'h21a30; force soc.dbg_do = 32'h41b785b3; #1000;
force soc.dbg_adr = 32'h21a34; force soc.dbg_do = 32'h2e070063; #1000;
force soc.dbg_adr = 32'h21a38; force soc.dbg_do = 32'h00bef463; #1000;
force soc.dbg_adr = 32'h21a3c; force soc.dbg_do = 32'h000e8593; #1000;
force soc.dbg_adr = 32'h21a40; force soc.dbg_do = 32'h0026f693; #1000;
force soc.dbg_adr = 32'h21a44; force soc.dbg_do = 32'h52068263; #1000;
force soc.dbg_adr = 32'h21a48; force soc.dbg_do = 32'h000c0713; #1000;
force soc.dbg_adr = 32'h21a4c; force soc.dbg_do = 32'h00200c93; #1000;
force soc.dbg_adr = 32'h21a50; force soc.dbg_do = 32'h03212023; #1000;
force soc.dbg_adr = 32'h21a54; force soc.dbg_do = 32'h03712423; #1000;
force soc.dbg_adr = 32'h21a58; force soc.dbg_do = 32'h00ee8c33; #1000;
force soc.dbg_adr = 32'h21a5c; force soc.dbg_do = 32'h01c12e23; #1000;
force soc.dbg_adr = 32'h21a60; force soc.dbg_do = 32'h03912223; #1000;
force soc.dbg_adr = 32'h21a64; force soc.dbg_do = 32'h00070793; #1000;
force soc.dbg_adr = 32'h21a68; force soc.dbg_do = 32'h01812b83; #1000;
force soc.dbg_adr = 32'h21a6c; force soc.dbg_do = 32'h00070913; #1000;
force soc.dbg_adr = 32'h21a70; force soc.dbg_do = 32'h00058d13; #1000;
force soc.dbg_adr = 32'h21a74; force soc.dbg_do = 32'h02fc0863; #1000;
force soc.dbg_adr = 32'h21a78; force soc.dbg_do = 32'h00048693; #1000;
force soc.dbg_adr = 32'h21a7c; force soc.dbg_do = 32'h00078613; #1000;
force soc.dbg_adr = 32'h21a80; force soc.dbg_do = 32'h000b8593; #1000;
force soc.dbg_adr = 32'h21a84; force soc.dbg_do = 32'h00178c93; #1000;
force soc.dbg_adr = 32'h21a88; force soc.dbg_do = 32'h000980e7; #1000;
force soc.dbg_adr = 32'h21a8c; force soc.dbg_do = 32'h412c8733; #1000;
force soc.dbg_adr = 32'h21a90; force soc.dbg_do = 32'h00ed8733; #1000;
force soc.dbg_adr = 32'h21a94; force soc.dbg_do = 32'h00074503; #1000;
force soc.dbg_adr = 32'h21a98; force soc.dbg_do = 32'h2e050e63; #1000;
force soc.dbg_adr = 32'h21a9c; force soc.dbg_do = 32'h000c8793; #1000;
force soc.dbg_adr = 32'h21aa0; force soc.dbg_do = 32'hfcfc1ce3; #1000;
force soc.dbg_adr = 32'h21aa4; force soc.dbg_do = 32'h01c12e03; #1000;
force soc.dbg_adr = 32'h21aa8; force soc.dbg_do = 32'h02012903; #1000;
force soc.dbg_adr = 32'h21aac; force soc.dbg_do = 32'h02412c83; #1000;
force soc.dbg_adr = 32'h21ab0; force soc.dbg_do = 32'h02812b83; #1000;
force soc.dbg_adr = 32'h21ab4; force soc.dbg_do = 32'h000d0593; #1000;
force soc.dbg_adr = 32'h21ab8; force soc.dbg_do = 32'h380c9263; #1000;
force soc.dbg_adr = 32'h21abc; force soc.dbg_do = 32'h07012d03; #1000;
force soc.dbg_adr = 32'h21ac0; force soc.dbg_do = 32'h00090d93; #1000;
force soc.dbg_adr = 32'h21ac4; force soc.dbg_do = 32'hba5ff06f; #1000;
force soc.dbg_adr = 32'h21ac8; force soc.dbg_do = 32'h0026f693; #1000;
force soc.dbg_adr = 32'h21acc; force soc.dbg_do = 32'h001c0c93; #1000;
force soc.dbg_adr = 32'h21ad0; force soc.dbg_do = 32'h004d8913; #1000;
force soc.dbg_adr = 32'h21ad4; force soc.dbg_do = 32'h2e068063; #1000;
force soc.dbg_adr = 32'h21ad8; force soc.dbg_do = 32'h000dc503; #1000;
force soc.dbg_adr = 32'h21adc; force soc.dbg_do = 32'h01812583; #1000;
force soc.dbg_adr = 32'h21ae0; force soc.dbg_do = 32'h01c12e23; #1000;
force soc.dbg_adr = 32'h21ae4; force soc.dbg_do = 32'h000c0613; #1000;
force soc.dbg_adr = 32'h21ae8; force soc.dbg_do = 32'h00048693; #1000;
force soc.dbg_adr = 32'h21aec; force soc.dbg_do = 32'h000980e7; #1000;
force soc.dbg_adr = 32'h21af0; force soc.dbg_do = 32'h01c12e03; #1000;
force soc.dbg_adr = 32'h21af4; force soc.dbg_do = 32'h00100793; #1000;
force soc.dbg_adr = 32'h21af8; force soc.dbg_do = 32'h01cc0c33; #1000;
force soc.dbg_adr = 32'h21afc; force soc.dbg_do = 32'h5bc7f263; #1000;
force soc.dbg_adr = 32'h21b00; force soc.dbg_do = 32'h07a12823; #1000;
force soc.dbg_adr = 32'h21b04; force soc.dbg_do = 32'h01812d03; #1000;
force soc.dbg_adr = 32'h21b08; force soc.dbg_do = 32'h000c8613; #1000;
force soc.dbg_adr = 32'h21b0c; force soc.dbg_do = 32'h00048693; #1000;
force soc.dbg_adr = 32'h21b10; force soc.dbg_do = 32'h001c8c93; #1000;
force soc.dbg_adr = 32'h21b14; force soc.dbg_do = 32'h000d0593; #1000;
force soc.dbg_adr = 32'h21b18; force soc.dbg_do = 32'h02000513; #1000;
force soc.dbg_adr = 32'h21b1c; force soc.dbg_do = 32'h000980e7; #1000;
force soc.dbg_adr = 32'h21b20; force soc.dbg_do = 32'hff8c94e3; #1000;
force soc.dbg_adr = 32'h21b24; force soc.dbg_do = 32'h07012d03; #1000;
force soc.dbg_adr = 32'h21b28; force soc.dbg_do = 32'h00090d93; #1000;
force soc.dbg_adr = 32'h21b2c; force soc.dbg_do = 32'hb3dff06f; #1000;
force soc.dbg_adr = 32'h21b30; force soc.dbg_do = 32'h07a12823; #1000;
force soc.dbg_adr = 32'h21b34; force soc.dbg_do = 32'h06f00793; #1000;
force soc.dbg_adr = 32'h21b38; force soc.dbg_do = 32'h32f50c63; #1000;
force soc.dbg_adr = 32'h21b3c; force soc.dbg_do = 32'h1aa7ea63; #1000;
force soc.dbg_adr = 32'h21b40; force soc.dbg_do = 32'h06900793; #1000;
force soc.dbg_adr = 32'h21b44; force soc.dbg_do = 32'hfef6f593; #1000;
force soc.dbg_adr = 32'h21b48; force soc.dbg_do = 32'h1af51ae3; #1000;
force soc.dbg_adr = 32'h21b4c; force soc.dbg_do = 32'h4006fd13; #1000;
force soc.dbg_adr = 32'h21b50; force soc.dbg_do = 32'h000d0663; #1000;
force soc.dbg_adr = 32'h21b54; force soc.dbg_do = 32'hfee6f593; #1000;
force soc.dbg_adr = 32'h21b58; force soc.dbg_do = 32'h40000d13; #1000;
force soc.dbg_adr = 32'h21b5c; force soc.dbg_do = 32'h2005f693; #1000;
force soc.dbg_adr = 32'h21b60; force soc.dbg_do = 32'h56069463; #1000;
force soc.dbg_adr = 32'h21b64; force soc.dbg_do = 32'h004d8793; #1000;
force soc.dbg_adr = 32'h21b68; force soc.dbg_do = 32'h1005fc93; #1000;
force soc.dbg_adr = 32'h21b6c; force soc.dbg_do = 32'h00f12e23; #1000;
force soc.dbg_adr = 32'h21b70; force soc.dbg_do = 32'h760c9e63; #1000;
force soc.dbg_adr = 32'h21b74; force soc.dbg_do = 32'h0405f713; #1000;
force soc.dbg_adr = 32'h21b78; force soc.dbg_do = 32'h74070863; #1000;
force soc.dbg_adr = 32'h21b7c; force soc.dbg_do = 32'h000dc703; #1000;
force soc.dbg_adr = 32'h21b80; force soc.dbg_do = 32'h00070693; #1000;
force soc.dbg_adr = 32'h21b84; force soc.dbg_do = 32'h01f75813; #1000;
force soc.dbg_adr = 32'h21b88; force soc.dbg_do = 32'h72070a63; #1000;
force soc.dbg_adr = 32'h21b8c; force soc.dbg_do = 32'h00068d13; #1000;
force soc.dbg_adr = 32'h21b90; force soc.dbg_do = 32'h04010713; #1000;
force soc.dbg_adr = 32'h21b94; force soc.dbg_do = 32'h03312623; #1000;
force soc.dbg_adr = 32'h21b98; force soc.dbg_do = 32'h02912823; #1000;
force soc.dbg_adr = 32'h21b9c; force soc.dbg_do = 32'h000c8993; #1000;
force soc.dbg_adr = 32'h21ba0; force soc.dbg_do = 32'h000d0493; #1000;
force soc.dbg_adr = 32'h21ba4; force soc.dbg_do = 32'h02000913; #1000;
force soc.dbg_adr = 32'h21ba8; force soc.dbg_do = 32'h03012023; #1000;
force soc.dbg_adr = 32'h21bac; force soc.dbg_do = 32'h03c12223; #1000;
force soc.dbg_adr = 32'h21bb0; force soc.dbg_do = 32'h03d12423; #1000;
force soc.dbg_adr = 32'h21bb4; force soc.dbg_do = 32'h00058d13; #1000;
force soc.dbg_adr = 32'h21bb8; force soc.dbg_do = 32'h000b8c93; #1000;
force soc.dbg_adr = 32'h21bbc; force soc.dbg_do = 32'h00070d93; #1000;
force soc.dbg_adr = 32'h21bc0; force soc.dbg_do = 32'h0080006f; #1000;
force soc.dbg_adr = 32'h21bc4; force soc.dbg_do = 32'h03298e63; #1000;
force soc.dbg_adr = 32'h21bc8; force soc.dbg_do = 32'h00a00593; #1000;
force soc.dbg_adr = 32'h21bcc; force soc.dbg_do = 32'h00048513; #1000;
force soc.dbg_adr = 32'h21bd0; force soc.dbg_do = 32'h6f5010ef; #1000;
force soc.dbg_adr = 32'h21bd4; force soc.dbg_do = 32'h00198993; #1000;
force soc.dbg_adr = 32'h21bd8; force soc.dbg_do = 32'h013d8bb3; #1000;
force soc.dbg_adr = 32'h21bdc; force soc.dbg_do = 32'h03050513; #1000;
force soc.dbg_adr = 32'h21be0; force soc.dbg_do = 32'hfeab8fa3; #1000;
force soc.dbg_adr = 32'h21be4; force soc.dbg_do = 32'h00a00593; #1000;
force soc.dbg_adr = 32'h21be8; force soc.dbg_do = 32'h00048513; #1000;
force soc.dbg_adr = 32'h21bec; force soc.dbg_do = 32'h691010ef; #1000;
force soc.dbg_adr = 32'h21bf0; force soc.dbg_do = 32'h00048b93; #1000;
force soc.dbg_adr = 32'h21bf4; force soc.dbg_do = 32'h00900793; #1000;
force soc.dbg_adr = 32'h21bf8; force soc.dbg_do = 32'h00050493; #1000;
force soc.dbg_adr = 32'h21bfc; force soc.dbg_do = 32'hfd77e4e3; #1000;
force soc.dbg_adr = 32'h21c00; force soc.dbg_do = 32'h000c8b93; #1000;
force soc.dbg_adr = 32'h21c04; force soc.dbg_do = 32'h02012803; #1000;
force soc.dbg_adr = 32'h21c08; force soc.dbg_do = 32'h00098c93; #1000;
force soc.dbg_adr = 32'h21c0c; force soc.dbg_do = 32'h02412e03; #1000;
force soc.dbg_adr = 32'h21c10; force soc.dbg_do = 32'h02812e83; #1000;
force soc.dbg_adr = 32'h21c14; force soc.dbg_do = 32'h03012483; #1000;
force soc.dbg_adr = 32'h21c18; force soc.dbg_do = 32'h02c12983; #1000;
force soc.dbg_adr = 32'h21c1c; force soc.dbg_do = 32'h000d0593; #1000;
force soc.dbg_adr = 32'h21c20; force soc.dbg_do = 32'h000d8713; #1000;
force soc.dbg_adr = 32'h21c24; force soc.dbg_do = 32'h00b12423; #1000;
force soc.dbg_adr = 32'h21c28; force soc.dbg_do = 32'h01c12223; #1000;
force soc.dbg_adr = 32'h21c2c; force soc.dbg_do = 32'h01d12023; #1000;
force soc.dbg_adr = 32'h21c30; force soc.dbg_do = 32'h000c8793; #1000;
force soc.dbg_adr = 32'h21c34; force soc.dbg_do = 32'h000c0613; #1000;
force soc.dbg_adr = 32'h21c38; force soc.dbg_do = 32'h00a00893; #1000;
force soc.dbg_adr = 32'h21c3c; force soc.dbg_do = 32'h01812583; #1000;
force soc.dbg_adr = 32'h21c40; force soc.dbg_do = 32'h00048693; #1000;
force soc.dbg_adr = 32'h21c44; force soc.dbg_do = 32'h00098513; #1000;
force soc.dbg_adr = 32'h21c48; force soc.dbg_do = 32'hc3cff0ef; #1000;
force soc.dbg_adr = 32'h21c4c; force soc.dbg_do = 32'h00050c13; #1000;
force soc.dbg_adr = 32'h21c50; force soc.dbg_do = 32'h01c12d83; #1000;
force soc.dbg_adr = 32'h21c54; force soc.dbg_do = 32'h07012d03; #1000;
force soc.dbg_adr = 32'h21c58; force soc.dbg_do = 32'ha11ff06f; #1000;
force soc.dbg_adr = 32'h21c5c; force soc.dbg_do = 32'h000c4503; #1000;
force soc.dbg_adr = 32'h21c60; force soc.dbg_do = 32'h000219b7; #1000;
force soc.dbg_adr = 32'h21c64; force soc.dbg_do = 32'h08098993; #1000;
force soc.dbg_adr = 32'h21c68; force soc.dbg_do = 32'h00000b93; #1000;
force soc.dbg_adr = 32'h21c6c; force soc.dbg_do = 32'h9a051ae3; #1000;
force soc.dbg_adr = 32'h21c70; force soc.dbg_do = 32'h00000413; #1000;
force soc.dbg_adr = 32'h21c74; force soc.dbg_do = 32'hc49be8e3; #1000;
force soc.dbg_adr = 32'h21c78; force soc.dbg_do = 32'hc49ff06f; #1000;
force soc.dbg_adr = 32'h21c7c; force soc.dbg_do = 32'h00078713; #1000;
force soc.dbg_adr = 32'h21c80; force soc.dbg_do = 32'h002e9793; #1000;
force soc.dbg_adr = 32'h21c84; force soc.dbg_do = 32'h01d787b3; #1000;
force soc.dbg_adr = 32'h21c88; force soc.dbg_do = 32'h00160613; #1000;
force soc.dbg_adr = 32'h21c8c; force soc.dbg_do = 32'h00179793; #1000;
force soc.dbg_adr = 32'h21c90; force soc.dbg_do = 32'h00a787b3; #1000;
force soc.dbg_adr = 32'h21c94; force soc.dbg_do = 32'h00064503; #1000;
force soc.dbg_adr = 32'h21c98; force soc.dbg_do = 32'hfd078e93; #1000;
force soc.dbg_adr = 32'h21c9c; force soc.dbg_do = 32'hfd050793; #1000;
force soc.dbg_adr = 32'h21ca0; force soc.dbg_do = 32'h0ff7f793; #1000;
force soc.dbg_adr = 32'h21ca4; force soc.dbg_do = 32'hfcf77ee3; #1000;
force soc.dbg_adr = 32'h21ca8; force soc.dbg_do = 32'h00060b93; #1000;
force soc.dbg_adr = 32'h21cac; force soc.dbg_do = 32'h00160713; #1000;
force soc.dbg_adr = 32'h21cb0; force soc.dbg_do = 32'ha19ff06f; #1000;
force soc.dbg_adr = 32'h21cb4; force soc.dbg_do = 32'h000dae83; #1000;
force soc.dbg_adr = 32'h21cb8; force soc.dbg_do = 32'h002bc503; #1000;
force soc.dbg_adr = 32'h21cbc; force soc.dbg_do = 32'h002b8b93; #1000;
force soc.dbg_adr = 32'h21cc0; force soc.dbg_do = 32'hfffec793; #1000;
force soc.dbg_adr = 32'h21cc4; force soc.dbg_do = 32'h41f7d793; #1000;
force soc.dbg_adr = 32'h21cc8; force soc.dbg_do = 32'h004d8d93; #1000;
force soc.dbg_adr = 32'h21ccc; force soc.dbg_do = 32'h00fefeb3; #1000;
force soc.dbg_adr = 32'h21cd0; force soc.dbg_do = 32'h001b8713; #1000;
force soc.dbg_adr = 32'h21cd4; force soc.dbg_do = 32'h9f5ff06f; #1000;
force soc.dbg_adr = 32'h21cd8; force soc.dbg_do = 32'hfef6f613; #1000;
force soc.dbg_adr = 32'h21cdc; force soc.dbg_do = 32'h4006f793; #1000;
force soc.dbg_adr = 32'h21ce0; force soc.dbg_do = 32'h02166613; #1000;
force soc.dbg_adr = 32'h21ce4; force soc.dbg_do = 32'h04010713; #1000;
force soc.dbg_adr = 32'h21ce8; force soc.dbg_do = 32'hb6079ee3; #1000;
force soc.dbg_adr = 32'h21cec; force soc.dbg_do = 32'hb39ff06f; #1000;
force soc.dbg_adr = 32'h21cf0; force soc.dbg_do = 32'h30c50863; #1000;
force soc.dbg_adr = 32'h21cf4; force soc.dbg_do = 32'h00a00613; #1000;
force soc.dbg_adr = 32'h21cf8; force soc.dbg_do = 32'hfef6f693; #1000;
force soc.dbg_adr = 32'h21cfc; force soc.dbg_do = 32'h00060893; #1000;
force soc.dbg_adr = 32'h21d00; force soc.dbg_do = 32'h00000f13; #1000;
force soc.dbg_adr = 32'h21d04; force soc.dbg_do = 32'ha79ff06f; #1000;
force soc.dbg_adr = 32'h21d08; force soc.dbg_do = 32'h4006f793; #1000;
force soc.dbg_adr = 32'h21d0c; force soc.dbg_do = 32'h41b605b3; #1000;
force soc.dbg_adr = 32'h21d10; force soc.dbg_do = 32'hd20794e3; #1000;
force soc.dbg_adr = 32'h21d14; force soc.dbg_do = 32'h0026f693; #1000;
force soc.dbg_adr = 32'h21d18; force soc.dbg_do = 32'h2c068863; #1000;
force soc.dbg_adr = 32'h21d1c; force soc.dbg_do = 32'h000c0713; #1000;
force soc.dbg_adr = 32'h21d20; force soc.dbg_do = 32'h00200c93; #1000;
force soc.dbg_adr = 32'h21d24; force soc.dbg_do = 32'h01812d03; #1000;
force soc.dbg_adr = 32'h21d28; force soc.dbg_do = 32'h000b8793; #1000;
force soc.dbg_adr = 32'h21d2c; force soc.dbg_do = 32'h03212023; #1000;
force soc.dbg_adr = 32'h21d30; force soc.dbg_do = 32'h01c12e23; #1000;
force soc.dbg_adr = 32'h21d34; force soc.dbg_do = 32'h00070913; #1000;
force soc.dbg_adr = 32'h21d38; force soc.dbg_do = 32'h02b12223; #1000;
force soc.dbg_adr = 32'h21d3c; force soc.dbg_do = 32'h00070b93; #1000;
force soc.dbg_adr = 32'h21d40; force soc.dbg_do = 32'h00078c13; #1000;
force soc.dbg_adr = 32'h21d44; force soc.dbg_do = 32'h000b8613; #1000;
force soc.dbg_adr = 32'h21d48; force soc.dbg_do = 32'h00048693; #1000;
force soc.dbg_adr = 32'h21d4c; force soc.dbg_do = 32'h000d0593; #1000;
force soc.dbg_adr = 32'h21d50; force soc.dbg_do = 32'h000980e7; #1000;
force soc.dbg_adr = 32'h21d54; force soc.dbg_do = 32'h001b8b93; #1000;
force soc.dbg_adr = 32'h21d58; force soc.dbg_do = 32'h412b8733; #1000;
force soc.dbg_adr = 32'h21d5c; force soc.dbg_do = 32'h00ed8733; #1000;
force soc.dbg_adr = 32'h21d60; force soc.dbg_do = 32'h00074503; #1000;
force soc.dbg_adr = 32'h21d64; force soc.dbg_do = 32'hfe0510e3; #1000;
force soc.dbg_adr = 32'h21d68; force soc.dbg_do = 32'h000c0793; #1000;
force soc.dbg_adr = 32'h21d6c; force soc.dbg_do = 32'h01c12e03; #1000;
force soc.dbg_adr = 32'h21d70; force soc.dbg_do = 32'h000b8c13; #1000;
force soc.dbg_adr = 32'h21d74; force soc.dbg_do = 32'h02012903; #1000;
force soc.dbg_adr = 32'h21d78; force soc.dbg_do = 32'h02412583; #1000;
force soc.dbg_adr = 32'h21d7c; force soc.dbg_do = 32'h00078b93; #1000;
force soc.dbg_adr = 32'h21d80; force soc.dbg_do = 32'hd39ff06f; #1000;
force soc.dbg_adr = 32'h21d84; force soc.dbg_do = 32'h002bc503; #1000;
force soc.dbg_adr = 32'h21d88; force soc.dbg_do = 32'h0c06e693; #1000;
force soc.dbg_adr = 32'h21d8c; force soc.dbg_do = 32'h003b8713; #1000;
force soc.dbg_adr = 32'h21d90; force soc.dbg_do = 32'h9a9ff06f; #1000;
force soc.dbg_adr = 32'h21d94; force soc.dbg_do = 32'h000d0593; #1000;
force soc.dbg_adr = 32'h21d98; force soc.dbg_do = 32'h000c8d13; #1000;
force soc.dbg_adr = 32'h21d9c; force soc.dbg_do = 32'h01c12e03; #1000;
force soc.dbg_adr = 32'h21da0; force soc.dbg_do = 32'h02012903; #1000;
force soc.dbg_adr = 32'h21da4; force soc.dbg_do = 32'h02412c83; #1000;
force soc.dbg_adr = 32'h21da8; force soc.dbg_do = 32'h02812b83; #1000;
force soc.dbg_adr = 32'h21dac; force soc.dbg_do = 32'h000d0c13; #1000;
force soc.dbg_adr = 32'h21db0; force soc.dbg_do = 32'hd09ff06f; #1000;
force soc.dbg_adr = 32'h21db4; force soc.dbg_do = 32'h00100793; #1000;
force soc.dbg_adr = 32'h21db8; force soc.dbg_do = 32'h2dc7fa63; #1000;
force soc.dbg_adr = 32'h21dbc; force soc.dbg_do = 32'h07a12823; #1000;
force soc.dbg_adr = 32'h21dc0; force soc.dbg_do = 32'h000b8d13; #1000;
force soc.dbg_adr = 32'h21dc4; force soc.dbg_do = 32'h01812b83; #1000;
force soc.dbg_adr = 32'h21dc8; force soc.dbg_do = 32'hfffc0793; #1000;
force soc.dbg_adr = 32'h21dcc; force soc.dbg_do = 32'h03212023; #1000;
force soc.dbg_adr = 32'h21dd0; force soc.dbg_do = 32'h01c78cb3; #1000;
force soc.dbg_adr = 32'h21dd4; force soc.dbg_do = 32'h01c12e23; #1000;
force soc.dbg_adr = 32'h21dd8; force soc.dbg_do = 32'h000c0913; #1000;
force soc.dbg_adr = 32'h21ddc; force soc.dbg_do = 32'h00090613; #1000;
force soc.dbg_adr = 32'h21de0; force soc.dbg_do = 32'h00048693; #1000;
force soc.dbg_adr = 32'h21de4; force soc.dbg_do = 32'h00190913; #1000;
force soc.dbg_adr = 32'h21de8; force soc.dbg_do = 32'h000b8593; #1000;
force soc.dbg_adr = 32'h21dec; force soc.dbg_do = 32'h02000513; #1000;
force soc.dbg_adr = 32'h21df0; force soc.dbg_do = 32'h000980e7; #1000;
force soc.dbg_adr = 32'h21df4; force soc.dbg_do = 32'hff9914e3; #1000;
force soc.dbg_adr = 32'h21df8; force soc.dbg_do = 32'h01c12e03; #1000;
force soc.dbg_adr = 32'h21dfc; force soc.dbg_do = 32'h000dc503; #1000;
force soc.dbg_adr = 32'h21e00; force soc.dbg_do = 32'h01812583; #1000;
force soc.dbg_adr = 32'h21e04; force soc.dbg_do = 32'h000d0b93; #1000;
force soc.dbg_adr = 32'h21e08; force soc.dbg_do = 32'h00090d13; #1000;
force soc.dbg_adr = 32'h21e0c; force soc.dbg_do = 32'h02012903; #1000;
force soc.dbg_adr = 32'h21e10; force soc.dbg_do = 32'h000d0613; #1000;
force soc.dbg_adr = 32'h21e14; force soc.dbg_do = 32'h00048693; #1000;
force soc.dbg_adr = 32'h21e18; force soc.dbg_do = 32'h01cc0c33; #1000;
force soc.dbg_adr = 32'h21e1c; force soc.dbg_do = 32'h00090d93; #1000;
force soc.dbg_adr = 32'h21e20; force soc.dbg_do = 32'h000980e7; #1000;
force soc.dbg_adr = 32'h21e24; force soc.dbg_do = 32'h07012d03; #1000;
force soc.dbg_adr = 32'h21e28; force soc.dbg_do = 32'h841ff06f; #1000;
force soc.dbg_adr = 32'h21e2c; force soc.dbg_do = 32'h4006f593; #1000;
force soc.dbg_adr = 32'h21e30; force soc.dbg_do = 32'h6a059c63; #1000;
force soc.dbg_adr = 32'h21e34; force soc.dbg_do = 32'h0026f693; #1000;
force soc.dbg_adr = 32'h21e38; force soc.dbg_do = 32'h1a068863; #1000;
force soc.dbg_adr = 32'h21e3c; force soc.dbg_do = 32'h000c0c93; #1000;
force soc.dbg_adr = 32'h21e40; force soc.dbg_do = 32'hc7c5fee3; #1000;
force soc.dbg_adr = 32'h21e44; force soc.dbg_do = 32'h01812d03; #1000;
force soc.dbg_adr = 32'h21e48; force soc.dbg_do = 32'h01cc0e33; #1000;
force soc.dbg_adr = 32'h21e4c; force soc.dbg_do = 32'h40be0c33; #1000;
force soc.dbg_adr = 32'h21e50; force soc.dbg_do = 32'h000c8613; #1000;
force soc.dbg_adr = 32'h21e54; force soc.dbg_do = 32'h00048693; #1000;
force soc.dbg_adr = 32'h21e58; force soc.dbg_do = 32'h001c8c93; #1000;
force soc.dbg_adr = 32'h21e5c; force soc.dbg_do = 32'h000d0593; #1000;
force soc.dbg_adr = 32'h21e60; force soc.dbg_do = 32'h02000513; #1000;
force soc.dbg_adr = 32'h21e64; force soc.dbg_do = 32'h000980e7; #1000;
force soc.dbg_adr = 32'h21e68; force soc.dbg_do = 32'hff8c94e3; #1000;
force soc.dbg_adr = 32'h21e6c; force soc.dbg_do = 32'hc51ff06f; #1000;
force soc.dbg_adr = 32'h21e70; force soc.dbg_do = 32'h00800613; #1000;
force soc.dbg_adr = 32'h21e74; force soc.dbg_do = 32'h00060893; #1000;
force soc.dbg_adr = 32'h21e78; force soc.dbg_do = 32'h00000f13; #1000;
force soc.dbg_adr = 32'h21e7c; force soc.dbg_do = 32'h901ff06f; #1000;
force soc.dbg_adr = 32'h21e80; force soc.dbg_do = 32'h00200613; #1000;
force soc.dbg_adr = 32'h21e84; force soc.dbg_do = 32'h07a12823; #1000;
force soc.dbg_adr = 32'h21e88; force soc.dbg_do = 32'h00060893; #1000;
force soc.dbg_adr = 32'h21e8c; force soc.dbg_do = 32'h00000f13; #1000;
force soc.dbg_adr = 32'h21e90; force soc.dbg_do = 32'h8edff06f; #1000;
force soc.dbg_adr = 32'h21e94; force soc.dbg_do = 32'h007d8d93; #1000;
force soc.dbg_adr = 32'h21e98; force soc.dbg_do = 32'hff8dfd93; #1000;
force soc.dbg_adr = 32'h21e9c; force soc.dbg_do = 32'h000daf83; #1000;
force soc.dbg_adr = 32'h21ea0; force soc.dbg_do = 32'h004dac83; #1000;
force soc.dbg_adr = 32'h21ea4; force soc.dbg_do = 32'h008d8d93; #1000;
force soc.dbg_adr = 32'h21ea8; force soc.dbg_do = 32'h019fe7b3; #1000;
force soc.dbg_adr = 32'h21eac; force soc.dbg_do = 32'h16078663; #1000;
force soc.dbg_adr = 32'h21eb0; force soc.dbg_do = 32'h00585713; #1000;
force soc.dbg_adr = 32'h21eb4; force soc.dbg_do = 32'h00177713; #1000;
force soc.dbg_adr = 32'h21eb8; force soc.dbg_do = 32'h06100793; #1000;
force soc.dbg_adr = 32'h21ebc; force soc.dbg_do = 32'h00070463; #1000;
force soc.dbg_adr = 32'h21ec0; force soc.dbg_do = 32'h04100793; #1000;
force soc.dbg_adr = 32'h21ec4; force soc.dbg_do = 32'hff678793; #1000;
force soc.dbg_adr = 32'h21ec8; force soc.dbg_do = 32'h04010713; #1000;
force soc.dbg_adr = 32'h21ecc; force soc.dbg_do = 32'h03812423; #1000;
force soc.dbg_adr = 32'h21ed0; force soc.dbg_do = 32'h03312823; #1000;
force soc.dbg_adr = 32'h21ed4; force soc.dbg_do = 32'h02912a23; #1000;
force soc.dbg_adr = 32'h21ed8; force soc.dbg_do = 32'h03712c23; #1000;
force soc.dbg_adr = 32'h21edc; force soc.dbg_do = 32'h03b12e23; #1000;
force soc.dbg_adr = 32'h21ee0; force soc.dbg_do = 32'h00000d13; #1000;
force soc.dbg_adr = 32'h21ee4; force soc.dbg_do = 32'h02000913; #1000;
force soc.dbg_adr = 32'h21ee8; force soc.dbg_do = 32'h01c12e23; #1000;
force soc.dbg_adr = 32'h21eec; force soc.dbg_do = 32'h03012023; #1000;
force soc.dbg_adr = 32'h21ef0; force soc.dbg_do = 32'h03d12223; #1000;
force soc.dbg_adr = 32'h21ef4; force soc.dbg_do = 32'h03112623; #1000;
force soc.dbg_adr = 32'h21ef8; force soc.dbg_do = 32'h000f8493; #1000;
force soc.dbg_adr = 32'h21efc; force soc.dbg_do = 32'h00060993; #1000;
force soc.dbg_adr = 32'h21f00; force soc.dbg_do = 32'h000f0c13; #1000;
force soc.dbg_adr = 32'h21f04; force soc.dbg_do = 32'h00070b93; #1000;
force soc.dbg_adr = 32'h21f08; force soc.dbg_do = 32'h00078d93; #1000;
force soc.dbg_adr = 32'h21f0c; force soc.dbg_do = 32'h00098613; #1000;
force soc.dbg_adr = 32'h21f10; force soc.dbg_do = 32'h00000693; #1000;
force soc.dbg_adr = 32'h21f14; force soc.dbg_do = 32'h00048513; #1000;
force soc.dbg_adr = 32'h21f18; force soc.dbg_do = 32'h000c8593; #1000;
force soc.dbg_adr = 32'h21f1c; force soc.dbg_do = 32'h571000ef; #1000;
force soc.dbg_adr = 32'h21f20; force soc.dbg_do = 32'h0ff57513; #1000;
force soc.dbg_adr = 32'h21f24; force soc.dbg_do = 32'h00900793; #1000;
force soc.dbg_adr = 32'h21f28; force soc.dbg_do = 32'h18a7ea63; #1000;
force soc.dbg_adr = 32'h21f2c; force soc.dbg_do = 32'h03050793; #1000;
force soc.dbg_adr = 32'h21f30; force soc.dbg_do = 32'h0ff7f793; #1000;
force soc.dbg_adr = 32'h21f34; force soc.dbg_do = 32'h001d0d13; #1000;
force soc.dbg_adr = 32'h21f38; force soc.dbg_do = 32'h01ab86b3; #1000;
force soc.dbg_adr = 32'h21f3c; force soc.dbg_do = 32'hfef68fa3; #1000;
force soc.dbg_adr = 32'h21f40; force soc.dbg_do = 32'h00098613; #1000;
force soc.dbg_adr = 32'h21f44; force soc.dbg_do = 32'h00000693; #1000;
force soc.dbg_adr = 32'h21f48; force soc.dbg_do = 32'h00048513; #1000;
force soc.dbg_adr = 32'h21f4c; force soc.dbg_do = 32'h000c8593; #1000;
force soc.dbg_adr = 32'h21f50; force soc.dbg_do = 32'h774000ef; #1000;
force soc.dbg_adr = 32'h21f54; force soc.dbg_do = 32'h119c0463; #1000;
force soc.dbg_adr = 32'h21f58; force soc.dbg_do = 32'h112d0463; #1000;
force soc.dbg_adr = 32'h21f5c; force soc.dbg_do = 32'h00050493; #1000;
force soc.dbg_adr = 32'h21f60; force soc.dbg_do = 32'h00058c93; #1000;
force soc.dbg_adr = 32'h21f64; force soc.dbg_do = 32'hfa9ff06f; #1000;
force soc.dbg_adr = 32'h21f68; force soc.dbg_do = 32'h40000d13; #1000;
force soc.dbg_adr = 32'h21f6c; force soc.dbg_do = 32'h15c5f063; #1000;
force soc.dbg_adr = 32'h21f70; force soc.dbg_do = 32'h018e0733; #1000;
force soc.dbg_adr = 32'h21f74; force soc.dbg_do = 32'h03712423; #1000;
force soc.dbg_adr = 32'h21f78; force soc.dbg_do = 32'h000c0b93; #1000;
force soc.dbg_adr = 32'h21f7c; force soc.dbg_do = 32'h01812c03; #1000;
force soc.dbg_adr = 32'h21f80; force soc.dbg_do = 32'h40b70733; #1000;
force soc.dbg_adr = 32'h21f84; force soc.dbg_do = 32'h03212223; #1000;
force soc.dbg_adr = 32'h21f88; force soc.dbg_do = 32'h01c12e23; #1000;
force soc.dbg_adr = 32'h21f8c; force soc.dbg_do = 32'h00048913; #1000;
force soc.dbg_adr = 32'h21f90; force soc.dbg_do = 32'h03d12023; #1000;
force soc.dbg_adr = 32'h21f94; force soc.dbg_do = 32'h00070493; #1000;
force soc.dbg_adr = 32'h21f98; force soc.dbg_do = 32'h000b8613; #1000;
force soc.dbg_adr = 32'h21f9c; force soc.dbg_do = 32'h00090693; #1000;
force soc.dbg_adr = 32'h21fa0; force soc.dbg_do = 32'h001b8b93; #1000;
force soc.dbg_adr = 32'h21fa4; force soc.dbg_do = 32'h000c0593; #1000;
force soc.dbg_adr = 32'h21fa8; force soc.dbg_do = 32'h02000513; #1000;
force soc.dbg_adr = 32'h21fac; force soc.dbg_do = 32'h000980e7; #1000;
force soc.dbg_adr = 32'h21fb0; force soc.dbg_do = 32'hfe9b94e3; #1000;
force soc.dbg_adr = 32'h21fb4; force soc.dbg_do = 32'h01c12e03; #1000;
force soc.dbg_adr = 32'h21fb8; force soc.dbg_do = 32'h000dc503; #1000;
force soc.dbg_adr = 32'h21fbc; force soc.dbg_do = 32'h00048713; #1000;
force soc.dbg_adr = 32'h21fc0; force soc.dbg_do = 32'h000b8c13; #1000;
force soc.dbg_adr = 32'h21fc4; force soc.dbg_do = 32'h00090493; #1000;
force soc.dbg_adr = 32'h21fc8; force soc.dbg_do = 32'h02012e83; #1000;
force soc.dbg_adr = 32'h21fcc; force soc.dbg_do = 32'h02412903; #1000;
force soc.dbg_adr = 32'h21fd0; force soc.dbg_do = 32'h02812b83; #1000;
force soc.dbg_adr = 32'h21fd4; force soc.dbg_do = 32'h001e0593; #1000;
force soc.dbg_adr = 32'h21fd8; force soc.dbg_do = 32'hae0502e3; #1000;
force soc.dbg_adr = 32'h21fdc; force soc.dbg_do = 32'ha60d1ae3; #1000;
force soc.dbg_adr = 32'h21fe0; force soc.dbg_do = 32'h00000c93; #1000;
force soc.dbg_adr = 32'h21fe4; force soc.dbg_do = 32'hd41ff06f; #1000;
force soc.dbg_adr = 32'h21fe8; force soc.dbg_do = 32'h00000d13; #1000;
force soc.dbg_adr = 32'h21fec; force soc.dbg_do = 32'hf9c5e2e3; #1000;
force soc.dbg_adr = 32'h21ff0; force soc.dbg_do = 32'h00158593; #1000;
force soc.dbg_adr = 32'h21ff4; force soc.dbg_do = 32'h000c0713; #1000;
force soc.dbg_adr = 32'h21ff8; force soc.dbg_do = 32'hd20516e3; #1000;
force soc.dbg_adr = 32'h21ffc; force soc.dbg_do = 32'hac1ff06f; #1000;
force soc.dbg_adr = 32'h22000; force soc.dbg_do = 32'h01000613; #1000;
force soc.dbg_adr = 32'h22004; force soc.dbg_do = 32'h00060893; #1000;
force soc.dbg_adr = 32'h22008; force soc.dbg_do = 32'h00000f13; #1000;
force soc.dbg_adr = 32'h2200c; force soc.dbg_do = 32'hf70ff06f; #1000;
force soc.dbg_adr = 32'h22010; force soc.dbg_do = 32'h000dcc83; #1000;
force soc.dbg_adr = 32'h22014; force soc.dbg_do = 32'hfa4ff06f; #1000;
force soc.dbg_adr = 32'h22018; force soc.dbg_do = 32'hfef87813; #1000;
force soc.dbg_adr = 32'h2201c; force soc.dbg_do = 32'he8058ae3; #1000;
force soc.dbg_adr = 32'h22020; force soc.dbg_do = 32'h00000d13; #1000;
force soc.dbg_adr = 32'h22024; force soc.dbg_do = 32'h04010713; #1000;
force soc.dbg_adr = 32'h22028; force soc.dbg_do = 32'h01012423; #1000;
force soc.dbg_adr = 32'h2202c; force soc.dbg_do = 32'h01c12223; #1000;
force soc.dbg_adr = 32'h22030; force soc.dbg_do = 32'h01d12023; #1000;
force soc.dbg_adr = 32'h22034; force soc.dbg_do = 32'h000d0793; #1000;
force soc.dbg_adr = 32'h22038; force soc.dbg_do = 32'h000c0613; #1000;
force soc.dbg_adr = 32'h2203c; force soc.dbg_do = 32'h00000813; #1000;
force soc.dbg_adr = 32'h22040; force soc.dbg_do = 32'h01812583; #1000;
force soc.dbg_adr = 32'h22044; force soc.dbg_do = 32'h00048693; #1000;
force soc.dbg_adr = 32'h22048; force soc.dbg_do = 32'h00098513; #1000;
force soc.dbg_adr = 32'h2204c; force soc.dbg_do = 32'h838ff0ef; #1000;
force soc.dbg_adr = 32'h22050; force soc.dbg_do = 32'h00050c13; #1000;
force soc.dbg_adr = 32'h22054; force soc.dbg_do = 32'h07012d03; #1000;
force soc.dbg_adr = 32'h22058; force soc.dbg_do = 32'he10ff06f; #1000;
force soc.dbg_adr = 32'h2205c; force soc.dbg_do = 32'hef34fee3; #1000;
force soc.dbg_adr = 32'h22060; force soc.dbg_do = 32'h000b8713; #1000;
force soc.dbg_adr = 32'h22064; force soc.dbg_do = 32'h01c12e03; #1000;
force soc.dbg_adr = 32'h22068; force soc.dbg_do = 32'h02012803; #1000;
force soc.dbg_adr = 32'h2206c; force soc.dbg_do = 32'h02412e83; #1000;
force soc.dbg_adr = 32'h22070; force soc.dbg_do = 32'h02812c03; #1000;
force soc.dbg_adr = 32'h22074; force soc.dbg_do = 32'h02c12883; #1000;
force soc.dbg_adr = 32'h22078; force soc.dbg_do = 32'h03012983; #1000;
force soc.dbg_adr = 32'h2207c; force soc.dbg_do = 32'h03412483; #1000;
force soc.dbg_adr = 32'h22080; force soc.dbg_do = 32'h03c12d83; #1000;
force soc.dbg_adr = 32'h22084; force soc.dbg_do = 32'h03812b83; #1000;
force soc.dbg_adr = 32'h22088; force soc.dbg_do = 32'hfa1ff06f; #1000;
force soc.dbg_adr = 32'h2208c; force soc.dbg_do = 32'h000dc503; #1000;
force soc.dbg_adr = 32'h22090; force soc.dbg_do = 32'h01812583; #1000;
force soc.dbg_adr = 32'h22094; force soc.dbg_do = 32'h000c0613; #1000;
force soc.dbg_adr = 32'h22098; force soc.dbg_do = 32'h00048693; #1000;
force soc.dbg_adr = 32'h2209c; force soc.dbg_do = 32'h000980e7; #1000;
force soc.dbg_adr = 32'h220a0; force soc.dbg_do = 32'h000c8c13; #1000;
force soc.dbg_adr = 32'h220a4; force soc.dbg_do = 32'h00090d93; #1000;
force soc.dbg_adr = 32'h220a8; force soc.dbg_do = 32'hdc0ff06f; #1000;
force soc.dbg_adr = 32'h220ac; force soc.dbg_do = 32'ha00508e3; #1000;
force soc.dbg_adr = 32'h220b0; force soc.dbg_do = 32'h00158593; #1000;
force soc.dbg_adr = 32'h220b4; force soc.dbg_do = 32'h000c0713; #1000;
force soc.dbg_adr = 32'h220b8; force soc.dbg_do = 32'h999ff06f; #1000;
force soc.dbg_adr = 32'h220bc; force soc.dbg_do = 32'h01b507b3; #1000;
force soc.dbg_adr = 32'h220c0; force soc.dbg_do = 32'h0ff7f793; #1000;
force soc.dbg_adr = 32'h220c4; force soc.dbg_do = 32'he71ff06f; #1000;
force soc.dbg_adr = 32'h220c8; force soc.dbg_do = 32'h007d8d93; #1000;
force soc.dbg_adr = 32'h220cc; force soc.dbg_do = 32'hff8dfd93; #1000;
force soc.dbg_adr = 32'h220d0; force soc.dbg_do = 32'h004da703; #1000;
force soc.dbg_adr = 32'h220d4; force soc.dbg_do = 32'h000da883; #1000;
force soc.dbg_adr = 32'h220d8; force soc.dbg_do = 32'h008d8d93; #1000;
force soc.dbg_adr = 32'h220dc; force soc.dbg_do = 32'h01f75913; #1000;
force soc.dbg_adr = 32'h220e0; force soc.dbg_do = 32'h00e8e7b3; #1000;
force soc.dbg_adr = 32'h220e4; force soc.dbg_do = 32'h3c078263; #1000;
force soc.dbg_adr = 32'h220e8; force soc.dbg_do = 32'h41f75793; #1000;
force soc.dbg_adr = 32'h220ec; force soc.dbg_do = 32'h0117c8b3; #1000;
force soc.dbg_adr = 32'h220f0; force soc.dbg_do = 32'h00e7cd33; #1000;
force soc.dbg_adr = 32'h220f4; force soc.dbg_do = 32'h40f88733; #1000;
force soc.dbg_adr = 32'h220f8; force soc.dbg_do = 32'h40fd07b3; #1000;
force soc.dbg_adr = 32'h220fc; force soc.dbg_do = 32'h00e8bd33; #1000;
force soc.dbg_adr = 32'h22100; force soc.dbg_do = 32'h41a78d33; #1000;
force soc.dbg_adr = 32'h22104; force soc.dbg_do = 32'h00070893; #1000;
force soc.dbg_adr = 32'h22108; force soc.dbg_do = 32'h00000c93; #1000;
force soc.dbg_adr = 32'h2210c; force soc.dbg_do = 32'h04010713; #1000;
force soc.dbg_adr = 32'h22110; force soc.dbg_do = 32'h03812623; #1000;
force soc.dbg_adr = 32'h22114; force soc.dbg_do = 32'h03312823; #1000;
force soc.dbg_adr = 32'h22118; force soc.dbg_do = 32'h02912a23; #1000;
force soc.dbg_adr = 32'h2211c; force soc.dbg_do = 32'h000d0c13; #1000;
force soc.dbg_adr = 32'h22120; force soc.dbg_do = 32'h01212e23; #1000;
force soc.dbg_adr = 32'h22124; force soc.dbg_do = 32'h000b8d13; #1000;
force soc.dbg_adr = 32'h22128; force soc.dbg_do = 32'h03c12023; #1000;
force soc.dbg_adr = 32'h2212c; force soc.dbg_do = 32'h02b12223; #1000;
force soc.dbg_adr = 32'h22130; force soc.dbg_do = 32'h03d12423; #1000;
force soc.dbg_adr = 32'h22134; force soc.dbg_do = 32'h000c8993; #1000;
force soc.dbg_adr = 32'h22138; force soc.dbg_do = 32'h00088b93; #1000;
force soc.dbg_adr = 32'h2213c; force soc.dbg_do = 32'h00070493; #1000;
force soc.dbg_adr = 32'h22140; force soc.dbg_do = 32'h00c0006f; #1000;
force soc.dbg_adr = 32'h22144; force soc.dbg_do = 32'h02000793; #1000;
force soc.dbg_adr = 32'h22148; force soc.dbg_do = 32'h04f98c63; #1000;
force soc.dbg_adr = 32'h2214c; force soc.dbg_do = 32'h00a00613; #1000;
force soc.dbg_adr = 32'h22150; force soc.dbg_do = 32'h00000693; #1000;
force soc.dbg_adr = 32'h22154; force soc.dbg_do = 32'h000b8513; #1000;
force soc.dbg_adr = 32'h22158; force soc.dbg_do = 32'h000c0593; #1000;
force soc.dbg_adr = 32'h2215c; force soc.dbg_do = 32'h331000ef; #1000;
force soc.dbg_adr = 32'h22160; force soc.dbg_do = 32'h00198993; #1000;
force soc.dbg_adr = 32'h22164; force soc.dbg_do = 32'h01348933; #1000;
force soc.dbg_adr = 32'h22168; force soc.dbg_do = 32'h03050513; #1000;
force soc.dbg_adr = 32'h2216c; force soc.dbg_do = 32'hfea90fa3; #1000;
force soc.dbg_adr = 32'h22170; force soc.dbg_do = 32'h000c0593; #1000;
force soc.dbg_adr = 32'h22174; force soc.dbg_do = 32'h000b8513; #1000;
force soc.dbg_adr = 32'h22178; force soc.dbg_do = 32'h00a00613; #1000;
force soc.dbg_adr = 32'h2217c; force soc.dbg_do = 32'h00000693; #1000;
force soc.dbg_adr = 32'h22180; force soc.dbg_do = 32'h544000ef; #1000;
force soc.dbg_adr = 32'h22184; force soc.dbg_do = 32'h000c0c93; #1000;
force soc.dbg_adr = 32'h22188; force soc.dbg_do = 32'h000b8913; #1000;
force soc.dbg_adr = 32'h2218c; force soc.dbg_do = 32'h00058c13; #1000;
force soc.dbg_adr = 32'h22190; force soc.dbg_do = 32'h00050b93; #1000;
force soc.dbg_adr = 32'h22194; force soc.dbg_do = 32'hfa0c98e3; #1000;
force soc.dbg_adr = 32'h22198; force soc.dbg_do = 32'h00900693; #1000;
force soc.dbg_adr = 32'h2219c; force soc.dbg_do = 32'hfb26e4e3; #1000;
force soc.dbg_adr = 32'h221a0; force soc.dbg_do = 32'h00098c93; #1000;
force soc.dbg_adr = 32'h221a4; force soc.dbg_do = 32'h00048713; #1000;
force soc.dbg_adr = 32'h221a8; force soc.dbg_do = 32'h01c12903; #1000;
force soc.dbg_adr = 32'h221ac; force soc.dbg_do = 32'h02012e03; #1000;
force soc.dbg_adr = 32'h221b0; force soc.dbg_do = 32'h02412583; #1000;
force soc.dbg_adr = 32'h221b4; force soc.dbg_do = 32'h02812e83; #1000;
force soc.dbg_adr = 32'h221b8; force soc.dbg_do = 32'h02c12c03; #1000;
force soc.dbg_adr = 32'h221bc; force soc.dbg_do = 32'h03012983; #1000;
force soc.dbg_adr = 32'h221c0; force soc.dbg_do = 32'h03412483; #1000;
force soc.dbg_adr = 32'h221c4; force soc.dbg_do = 32'h000d0b93; #1000;
force soc.dbg_adr = 32'h221c8; force soc.dbg_do = 32'h00b12423; #1000;
force soc.dbg_adr = 32'h221cc; force soc.dbg_do = 32'h01c12223; #1000;
force soc.dbg_adr = 32'h221d0; force soc.dbg_do = 32'h01d12023; #1000;
force soc.dbg_adr = 32'h221d4; force soc.dbg_do = 32'h00090813; #1000;
force soc.dbg_adr = 32'h221d8; force soc.dbg_do = 32'h000c8793; #1000;
force soc.dbg_adr = 32'h221dc; force soc.dbg_do = 32'h000c0613; #1000;
force soc.dbg_adr = 32'h221e0; force soc.dbg_do = 32'h00a00893; #1000;
force soc.dbg_adr = 32'h221e4; force soc.dbg_do = 32'he5dff06f; #1000;
force soc.dbg_adr = 32'h221e8; force soc.dbg_do = 32'h00585713; #1000;
force soc.dbg_adr = 32'h221ec; force soc.dbg_do = 32'h00177713; #1000;
force soc.dbg_adr = 32'h221f0; force soc.dbg_do = 32'h06100793; #1000;
force soc.dbg_adr = 32'h221f4; force soc.dbg_do = 32'h00070463; #1000;
force soc.dbg_adr = 32'h221f8; force soc.dbg_do = 32'h04100793; #1000;
force soc.dbg_adr = 32'h221fc; force soc.dbg_do = 32'h000b8693; #1000;
force soc.dbg_adr = 32'h22200; force soc.dbg_do = 32'hff678793; #1000;
force soc.dbg_adr = 32'h22204; force soc.dbg_do = 32'h04010713; #1000;
force soc.dbg_adr = 32'h22208; force soc.dbg_do = 32'h03812623; #1000;
force soc.dbg_adr = 32'h2220c; force soc.dbg_do = 32'h03312823; #1000;
force soc.dbg_adr = 32'h22210; force soc.dbg_do = 32'h02912a23; #1000;
force soc.dbg_adr = 32'h22214; force soc.dbg_do = 32'h000d0b93; #1000;
force soc.dbg_adr = 32'h22218; force soc.dbg_do = 32'h00900d93; #1000;
force soc.dbg_adr = 32'h2221c; force soc.dbg_do = 32'h02000913; #1000;
force soc.dbg_adr = 32'h22220; force soc.dbg_do = 32'h03c12023; #1000;
force soc.dbg_adr = 32'h22224; force soc.dbg_do = 32'h03012223; #1000;
force soc.dbg_adr = 32'h22228; force soc.dbg_do = 32'h03d12423; #1000;
force soc.dbg_adr = 32'h2222c; force soc.dbg_do = 32'h00088993; #1000;
force soc.dbg_adr = 32'h22230; force soc.dbg_do = 32'h00070c13; #1000;
force soc.dbg_adr = 32'h22234; force soc.dbg_do = 32'h00078493; #1000;
force soc.dbg_adr = 32'h22238; force soc.dbg_do = 32'h00068d13; #1000;
force soc.dbg_adr = 32'h2223c; force soc.dbg_do = 32'h0300006f; #1000;
force soc.dbg_adr = 32'h22240; force soc.dbg_do = 32'h03078793; #1000;
force soc.dbg_adr = 32'h22244; force soc.dbg_do = 32'h0ff7f793; #1000;
force soc.dbg_adr = 32'h22248; force soc.dbg_do = 32'h001b8b93; #1000;
force soc.dbg_adr = 32'h2224c; force soc.dbg_do = 32'h017c06b3; #1000;
force soc.dbg_adr = 32'h22250; force soc.dbg_do = 32'hfef68fa3; #1000;
force soc.dbg_adr = 32'h22254; force soc.dbg_do = 32'h00098593; #1000;
force soc.dbg_adr = 32'h22258; force soc.dbg_do = 32'h000c8513; #1000;
force soc.dbg_adr = 32'h2225c; force soc.dbg_do = 32'h021010ef; #1000;
force soc.dbg_adr = 32'h22260; force soc.dbg_do = 32'h033ce663; #1000;
force soc.dbg_adr = 32'h22264; force soc.dbg_do = 32'h032b8463; #1000;
force soc.dbg_adr = 32'h22268; force soc.dbg_do = 32'h00050c93; #1000;
force soc.dbg_adr = 32'h2226c; force soc.dbg_do = 32'h00098593; #1000;
force soc.dbg_adr = 32'h22270; force soc.dbg_do = 32'h000c8513; #1000;
force soc.dbg_adr = 32'h22274; force soc.dbg_do = 32'h051010ef; #1000;
force soc.dbg_adr = 32'h22278; force soc.dbg_do = 32'h0ff57793; #1000;
force soc.dbg_adr = 32'h2227c; force soc.dbg_do = 32'hfcadf2e3; #1000;
force soc.dbg_adr = 32'h22280; force soc.dbg_do = 32'h009787b3; #1000;
force soc.dbg_adr = 32'h22284; force soc.dbg_do = 32'h0ff7f793; #1000;
force soc.dbg_adr = 32'h22288; force soc.dbg_do = 32'hfc1ff06f; #1000;
force soc.dbg_adr = 32'h2228c; force soc.dbg_do = 32'h000d0793; #1000;
force soc.dbg_adr = 32'h22290; force soc.dbg_do = 32'h00098893; #1000;
force soc.dbg_adr = 32'h22294; force soc.dbg_do = 32'h000b8d13; #1000;
force soc.dbg_adr = 32'h22298; force soc.dbg_do = 32'h000c0713; #1000;
force soc.dbg_adr = 32'h2229c; force soc.dbg_do = 32'h02012e03; #1000;
force soc.dbg_adr = 32'h222a0; force soc.dbg_do = 32'h02412803; #1000;
force soc.dbg_adr = 32'h222a4; force soc.dbg_do = 32'h02812e83; #1000;
force soc.dbg_adr = 32'h222a8; force soc.dbg_do = 32'h03012983; #1000;
force soc.dbg_adr = 32'h222ac; force soc.dbg_do = 32'h03412483; #1000;
force soc.dbg_adr = 32'h222b0; force soc.dbg_do = 32'h02c12c03; #1000;
force soc.dbg_adr = 32'h222b4; force soc.dbg_do = 32'h00078b93; #1000;
force soc.dbg_adr = 32'h222b8; force soc.dbg_do = 32'hd14ff06f; #1000;
force soc.dbg_adr = 32'h222bc; force soc.dbg_do = 32'h04010713; #1000;
force soc.dbg_adr = 32'h222c0; force soc.dbg_do = 32'h960d12e3; #1000;
force soc.dbg_adr = 32'h222c4; force soc.dbg_do = 32'h8cdff06f; #1000;
force soc.dbg_adr = 32'h222c8; force soc.dbg_do = 32'h0805f713; #1000;
force soc.dbg_adr = 32'h222cc; force soc.dbg_do = 32'h1e070463; #1000;
force soc.dbg_adr = 32'h222d0; force soc.dbg_do = 32'h000d9703; #1000;
force soc.dbg_adr = 32'h222d4; force soc.dbg_do = 32'h40f75513; #1000;
force soc.dbg_adr = 32'h222d8; force soc.dbg_do = 32'h00a746b3; #1000;
force soc.dbg_adr = 32'h222dc; force soc.dbg_do = 32'h40a686b3; #1000;
force soc.dbg_adr = 32'h222e0; force soc.dbg_do = 32'h01069693; #1000;
force soc.dbg_adr = 32'h222e4; force soc.dbg_do = 32'h0106d693; #1000;
force soc.dbg_adr = 32'h222e8; force soc.dbg_do = 32'h89dff06f; #1000;
force soc.dbg_adr = 32'h222ec; force soc.dbg_do = 32'h000da783; #1000;
force soc.dbg_adr = 32'h222f0; force soc.dbg_do = 32'h01f7d913; #1000;
force soc.dbg_adr = 32'h222f4; force soc.dbg_do = 32'h1c078a63; #1000;
force soc.dbg_adr = 32'h222f8; force soc.dbg_do = 32'h41f7d713; #1000;
force soc.dbg_adr = 32'h222fc; force soc.dbg_do = 32'h00f74d33; #1000;
force soc.dbg_adr = 32'h22300; force soc.dbg_do = 32'h40ed0d33; #1000;
force soc.dbg_adr = 32'h22304; force soc.dbg_do = 32'h04010713; #1000;
force soc.dbg_adr = 32'h22308; force soc.dbg_do = 32'h03212023; #1000;
force soc.dbg_adr = 32'h2230c; force soc.dbg_do = 32'h00900c93; #1000;
force soc.dbg_adr = 32'h22310; force soc.dbg_do = 32'h000d0913; #1000;
force soc.dbg_adr = 32'h22314; force soc.dbg_do = 32'h03c12223; #1000;
force soc.dbg_adr = 32'h22318; force soc.dbg_do = 32'h000b8d13; #1000;
force soc.dbg_adr = 32'h2231c; force soc.dbg_do = 32'h02b12423; #1000;
force soc.dbg_adr = 32'h22320; force soc.dbg_do = 32'h00048b93; #1000;
force soc.dbg_adr = 32'h22324; force soc.dbg_do = 32'h03d12623; #1000;
force soc.dbg_adr = 32'h22328; force soc.dbg_do = 32'h03312823; #1000;
force soc.dbg_adr = 32'h2232c; force soc.dbg_do = 32'h00068493; #1000;
force soc.dbg_adr = 32'h22330; force soc.dbg_do = 32'h00070d93; #1000;
force soc.dbg_adr = 32'h22334; force soc.dbg_do = 32'h00c0006f; #1000;
force soc.dbg_adr = 32'h22338; force soc.dbg_do = 32'h02000793; #1000;
force soc.dbg_adr = 32'h2233c; force soc.dbg_do = 32'h02f48c63; #1000;
force soc.dbg_adr = 32'h22340; force soc.dbg_do = 32'h00a00593; #1000;
force soc.dbg_adr = 32'h22344; force soc.dbg_do = 32'h00090513; #1000;
force soc.dbg_adr = 32'h22348; force soc.dbg_do = 32'h77c010ef; #1000;
force soc.dbg_adr = 32'h2234c; force soc.dbg_do = 32'h00148493; #1000;
force soc.dbg_adr = 32'h22350; force soc.dbg_do = 32'h009d89b3; #1000;
force soc.dbg_adr = 32'h22354; force soc.dbg_do = 32'h03050513; #1000;
force soc.dbg_adr = 32'h22358; force soc.dbg_do = 32'hfea98fa3; #1000;
force soc.dbg_adr = 32'h2235c; force soc.dbg_do = 32'h00a00593; #1000;
force soc.dbg_adr = 32'h22360; force soc.dbg_do = 32'h00090513; #1000;
force soc.dbg_adr = 32'h22364; force soc.dbg_do = 32'h00090993; #1000;
force soc.dbg_adr = 32'h22368; force soc.dbg_do = 32'h714010ef; #1000;
force soc.dbg_adr = 32'h2236c; force soc.dbg_do = 32'h00050913; #1000;
force soc.dbg_adr = 32'h22370; force soc.dbg_do = 32'hfd3ce4e3; #1000;
force soc.dbg_adr = 32'h22374; force soc.dbg_do = 32'h02012903; #1000;
force soc.dbg_adr = 32'h22378; force soc.dbg_do = 32'h02412e03; #1000;
force soc.dbg_adr = 32'h2237c; force soc.dbg_do = 32'h02812583; #1000;
force soc.dbg_adr = 32'h22380; force soc.dbg_do = 32'h02c12e83; #1000;
force soc.dbg_adr = 32'h22384; force soc.dbg_do = 32'h03012983; #1000;
force soc.dbg_adr = 32'h22388; force soc.dbg_do = 32'h00048693; #1000;
force soc.dbg_adr = 32'h2238c; force soc.dbg_do = 32'h000d8713; #1000;
force soc.dbg_adr = 32'h22390; force soc.dbg_do = 32'h000b8493; #1000;
force soc.dbg_adr = 32'h22394; force soc.dbg_do = 32'h000d0b93; #1000;
force soc.dbg_adr = 32'h22398; force soc.dbg_do = 32'h00b12423; #1000;
force soc.dbg_adr = 32'h2239c; force soc.dbg_do = 32'h01c12223; #1000;
force soc.dbg_adr = 32'h223a0; force soc.dbg_do = 32'h01d12023; #1000;
force soc.dbg_adr = 32'h223a4; force soc.dbg_do = 32'h00090813; #1000;
force soc.dbg_adr = 32'h223a8; force soc.dbg_do = 32'h00068793; #1000;
force soc.dbg_adr = 32'h223ac; force soc.dbg_do = 32'h000c0613; #1000;
force soc.dbg_adr = 32'h223b0; force soc.dbg_do = 32'h00a00893; #1000;
force soc.dbg_adr = 32'h223b4; force soc.dbg_do = 32'h889ff06f; #1000;
force soc.dbg_adr = 32'h223b8; force soc.dbg_do = 32'h000dad83; #1000;
force soc.dbg_adr = 32'h223bc; force soc.dbg_do = 32'h000d9863; #1000;
force soc.dbg_adr = 32'h223c0; force soc.dbg_do = 32'hfef87813; #1000;
force soc.dbg_adr = 32'h223c4; force soc.dbg_do = 32'h04010713; #1000;
force soc.dbg_adr = 32'h223c8; force soc.dbg_do = 32'h0c059663; #1000;
force soc.dbg_adr = 32'h223cc; force soc.dbg_do = 32'h00585693; #1000;
force soc.dbg_adr = 32'h223d0; force soc.dbg_do = 32'h0016f693; #1000;
force soc.dbg_adr = 32'h223d4; force soc.dbg_do = 32'h06100713; #1000;
force soc.dbg_adr = 32'h223d8; force soc.dbg_do = 32'h00068463; #1000;
force soc.dbg_adr = 32'h223dc; force soc.dbg_do = 32'h04100713; #1000;
force soc.dbg_adr = 32'h223e0; force soc.dbg_do = 32'hff670793; #1000;
force soc.dbg_adr = 32'h223e4; force soc.dbg_do = 32'h04010713; #1000;
force soc.dbg_adr = 32'h223e8; force soc.dbg_do = 32'h03812623; #1000;
force soc.dbg_adr = 32'h223ec; force soc.dbg_do = 32'h03312823; #1000;
force soc.dbg_adr = 32'h223f0; force soc.dbg_do = 32'h02912a23; #1000;
force soc.dbg_adr = 32'h223f4; force soc.dbg_do = 32'h000c8993; #1000;
force soc.dbg_adr = 32'h223f8; force soc.dbg_do = 32'h00900d13; #1000;
force soc.dbg_adr = 32'h223fc; force soc.dbg_do = 32'h000b8c93; #1000;
force soc.dbg_adr = 32'h22400; force soc.dbg_do = 32'h02000913; #1000;
force soc.dbg_adr = 32'h22404; force soc.dbg_do = 32'h03c12023; #1000;
force soc.dbg_adr = 32'h22408; force soc.dbg_do = 32'h03012223; #1000;
force soc.dbg_adr = 32'h2240c; force soc.dbg_do = 32'h03d12423; #1000;
force soc.dbg_adr = 32'h22410; force soc.dbg_do = 32'h00088c13; #1000;
force soc.dbg_adr = 32'h22414; force soc.dbg_do = 32'h00070493; #1000;
force soc.dbg_adr = 32'h22418; force soc.dbg_do = 32'h00078b93; #1000;
force soc.dbg_adr = 32'h2241c; force soc.dbg_do = 32'h0300006f; #1000;
force soc.dbg_adr = 32'h22420; force soc.dbg_do = 32'h03078793; #1000;
force soc.dbg_adr = 32'h22424; force soc.dbg_do = 32'h0ff7f793; #1000;
force soc.dbg_adr = 32'h22428; force soc.dbg_do = 32'h00198993; #1000;
force soc.dbg_adr = 32'h2242c; force soc.dbg_do = 32'h013486b3; #1000;
force soc.dbg_adr = 32'h22430; force soc.dbg_do = 32'hfef68fa3; #1000;
force soc.dbg_adr = 32'h22434; force soc.dbg_do = 32'h000c0593; #1000;
force soc.dbg_adr = 32'h22438; force soc.dbg_do = 32'h000d8513; #1000;
force soc.dbg_adr = 32'h2243c; force soc.dbg_do = 32'h640010ef; #1000;
force soc.dbg_adr = 32'h22440; force soc.dbg_do = 32'h038de663; #1000;
force soc.dbg_adr = 32'h22444; force soc.dbg_do = 32'h03298463; #1000;
force soc.dbg_adr = 32'h22448; force soc.dbg_do = 32'h00050d93; #1000;
force soc.dbg_adr = 32'h2244c; force soc.dbg_do = 32'h000c0593; #1000;
force soc.dbg_adr = 32'h22450; force soc.dbg_do = 32'h000d8513; #1000;
force soc.dbg_adr = 32'h22454; force soc.dbg_do = 32'h670010ef; #1000;
force soc.dbg_adr = 32'h22458; force soc.dbg_do = 32'h0ff57793; #1000;
force soc.dbg_adr = 32'h2245c; force soc.dbg_do = 32'hfcad72e3; #1000;
force soc.dbg_adr = 32'h22460; force soc.dbg_do = 32'h017787b3; #1000;
force soc.dbg_adr = 32'h22464; force soc.dbg_do = 32'h0ff7f793; #1000;
force soc.dbg_adr = 32'h22468; force soc.dbg_do = 32'hfc1ff06f; #1000;
force soc.dbg_adr = 32'h2246c; force soc.dbg_do = 32'h000c0893; #1000;
force soc.dbg_adr = 32'h22470; force soc.dbg_do = 32'h000c8b93; #1000;
force soc.dbg_adr = 32'h22474; force soc.dbg_do = 32'h00048713; #1000;
force soc.dbg_adr = 32'h22478; force soc.dbg_do = 32'h00098c93; #1000;
force soc.dbg_adr = 32'h2247c; force soc.dbg_do = 32'h02012e03; #1000;
force soc.dbg_adr = 32'h22480; force soc.dbg_do = 32'h02412803; #1000;
force soc.dbg_adr = 32'h22484; force soc.dbg_do = 32'h02812e83; #1000;
force soc.dbg_adr = 32'h22488; force soc.dbg_do = 32'h02c12c03; #1000;
force soc.dbg_adr = 32'h2248c; force soc.dbg_do = 32'h03012983; #1000;
force soc.dbg_adr = 32'h22490; force soc.dbg_do = 32'h03412483; #1000;
force soc.dbg_adr = 32'h22494; force soc.dbg_do = 32'h01012423; #1000;
force soc.dbg_adr = 32'h22498; force soc.dbg_do = 32'h01c12223; #1000;
force soc.dbg_adr = 32'h2249c; force soc.dbg_do = 32'h01d12023; #1000;
force soc.dbg_adr = 32'h224a0; force soc.dbg_do = 32'h000c8793; #1000;
force soc.dbg_adr = 32'h224a4; force soc.dbg_do = 32'hb38ff06f; #1000;
force soc.dbg_adr = 32'h224a8; force soc.dbg_do = 32'h020d1a63; #1000;
force soc.dbg_adr = 32'h224ac; force soc.dbg_do = 32'h00000893; #1000;
force soc.dbg_adr = 32'h224b0; force soc.dbg_do = 32'hc59ff06f; #1000;
force soc.dbg_adr = 32'h224b4; force soc.dbg_do = 32'h000da703; #1000;
force soc.dbg_adr = 32'h224b8; force soc.dbg_do = 32'h41f75513; #1000;
force soc.dbg_adr = 32'h224bc; force soc.dbg_do = 32'h00e546b3; #1000;
force soc.dbg_adr = 32'h224c0; force soc.dbg_do = 32'h40a686b3; #1000;
force soc.dbg_adr = 32'h224c4; force soc.dbg_do = 32'hec0ff06f; #1000;
force soc.dbg_adr = 32'h224c8; force soc.dbg_do = 32'h04010713; #1000;
force soc.dbg_adr = 32'h224cc; force soc.dbg_do = 32'hec0d16e3; #1000;
force soc.dbg_adr = 32'h224d0; force soc.dbg_do = 32'he35ff06f; #1000;
force soc.dbg_adr = 32'h224d4; force soc.dbg_do = 32'h000dac83; #1000;
force soc.dbg_adr = 32'h224d8; force soc.dbg_do = 32'hae0ff06f; #1000;
force soc.dbg_adr = 32'h224dc; force soc.dbg_do = 32'h00000c93; #1000;
force soc.dbg_adr = 32'h224e0; force soc.dbg_do = 32'h04010713; #1000;
force soc.dbg_adr = 32'h224e4; force soc.dbg_do = 32'hce5ff06f; #1000;
force soc.dbg_adr = 32'h224e8; force soc.dbg_do = 32'h0026f593; #1000;
force soc.dbg_adr = 32'h224ec; force soc.dbg_do = 32'ha6058ee3; #1000;
force soc.dbg_adr = 32'h224f0; force soc.dbg_do = 32'h000c0c93; #1000;
force soc.dbg_adr = 32'h224f4; force soc.dbg_do = 32'h00000593; #1000;
force soc.dbg_adr = 32'h224f8; force soc.dbg_do = 32'h949ff06f; #1000;
force soc.dbg_adr = 32'h224fc; force soc.dbg_do = 32'h06400793; #1000;
force soc.dbg_adr = 32'h22500; force soc.dbg_do = 32'he4f50663; #1000;
force soc.dbg_adr = 32'h22504; force soc.dbg_do = 32'h00a00613; #1000;
force soc.dbg_adr = 32'h22508; force soc.dbg_do = 32'h00058693; #1000;
force soc.dbg_adr = 32'h2250c; force soc.dbg_do = 32'h00060893; #1000;
force soc.dbg_adr = 32'h22510; force soc.dbg_do = 32'h00000f13; #1000;
force soc.dbg_adr = 32'h22514; force soc.dbg_do = 32'ha68ff06f; #1000;
force soc.dbg_adr = 32'h22518; force soc.dbg_do = 32'hfc010113; #1000;
force soc.dbg_adr = 32'h2251c; force soc.dbg_do = 32'h02410313; #1000;
force soc.dbg_adr = 32'h22520; force soc.dbg_do = 32'h00021e37; #1000;
force soc.dbg_adr = 32'h22524; force soc.dbg_do = 32'h02b12223; #1000;
force soc.dbg_adr = 32'h22528; force soc.dbg_do = 32'h02c12423; #1000;
force soc.dbg_adr = 32'h2252c; force soc.dbg_do = 32'h02d12623; #1000;
force soc.dbg_adr = 32'h22530; force soc.dbg_do = 32'h02e12823; #1000;
force soc.dbg_adr = 32'h22534; force soc.dbg_do = 32'h00050693; #1000;
force soc.dbg_adr = 32'h22538; force soc.dbg_do = 32'h00810593; #1000;
force soc.dbg_adr = 32'h2253c; force soc.dbg_do = 32'h00030713; #1000;
force soc.dbg_adr = 32'h22540; force soc.dbg_do = 32'h5bce0513; #1000;
force soc.dbg_adr = 32'h22544; force soc.dbg_do = 32'hfff00613; #1000;
force soc.dbg_adr = 32'h22548; force soc.dbg_do = 32'h00112e23; #1000;
force soc.dbg_adr = 32'h2254c; force soc.dbg_do = 32'h02f12a23; #1000;
force soc.dbg_adr = 32'h22550; force soc.dbg_do = 32'h03012c23; #1000;
force soc.dbg_adr = 32'h22554; force soc.dbg_do = 32'h03112e23; #1000;
force soc.dbg_adr = 32'h22558; force soc.dbg_do = 32'h00612623; #1000;
force soc.dbg_adr = 32'h2255c; force soc.dbg_do = 32'h880ff0ef; #1000;
force soc.dbg_adr = 32'h22560; force soc.dbg_do = 32'h01c12083; #1000;
force soc.dbg_adr = 32'h22564; force soc.dbg_do = 32'h04010113; #1000;
force soc.dbg_adr = 32'h22568; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h2256c; force soc.dbg_do = 32'hfc010113; #1000;
force soc.dbg_adr = 32'h22570; force soc.dbg_do = 32'h02810313; #1000;
force soc.dbg_adr = 32'h22574; force soc.dbg_do = 32'h00058e93; #1000;
force soc.dbg_adr = 32'h22578; force soc.dbg_do = 32'h00021e37; #1000;
force soc.dbg_adr = 32'h2257c; force soc.dbg_do = 32'h02c12423; #1000;
force soc.dbg_adr = 32'h22580; force soc.dbg_do = 32'h02d12623; #1000;
force soc.dbg_adr = 32'h22584; force soc.dbg_do = 32'h02e12823; #1000;
force soc.dbg_adr = 32'h22588; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h2258c; force soc.dbg_do = 32'h000e8693; #1000;
force soc.dbg_adr = 32'h22590; force soc.dbg_do = 32'h00030713; #1000;
force soc.dbg_adr = 32'h22594; force soc.dbg_do = 32'h070e0513; #1000;
force soc.dbg_adr = 32'h22598; force soc.dbg_do = 32'hfff00613; #1000;
force soc.dbg_adr = 32'h2259c; force soc.dbg_do = 32'h00112e23; #1000;
force soc.dbg_adr = 32'h225a0; force soc.dbg_do = 32'h02f12a23; #1000;
force soc.dbg_adr = 32'h225a4; force soc.dbg_do = 32'h03012c23; #1000;
force soc.dbg_adr = 32'h225a8; force soc.dbg_do = 32'h03112e23; #1000;
force soc.dbg_adr = 32'h225ac; force soc.dbg_do = 32'h00612623; #1000;
force soc.dbg_adr = 32'h225b0; force soc.dbg_do = 32'h82cff0ef; #1000;
force soc.dbg_adr = 32'h225b4; force soc.dbg_do = 32'h01c12083; #1000;
force soc.dbg_adr = 32'h225b8; force soc.dbg_do = 32'h04010113; #1000;
force soc.dbg_adr = 32'h225bc; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h225c0; force soc.dbg_do = 32'hfc010113; #1000;
force soc.dbg_adr = 32'h225c4; force soc.dbg_do = 32'h02c10313; #1000;
force soc.dbg_adr = 32'h225c8; force soc.dbg_do = 32'h00058f13; #1000;
force soc.dbg_adr = 32'h225cc; force soc.dbg_do = 32'h00060e93; #1000;
force soc.dbg_adr = 32'h225d0; force soc.dbg_do = 32'h00021e37; #1000;
force soc.dbg_adr = 32'h225d4; force soc.dbg_do = 32'h02d12623; #1000;
force soc.dbg_adr = 32'h225d8; force soc.dbg_do = 32'h02e12823; #1000;
force soc.dbg_adr = 32'h225dc; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h225e0; force soc.dbg_do = 32'h000f0613; #1000;
force soc.dbg_adr = 32'h225e4; force soc.dbg_do = 32'h000e8693; #1000;
force soc.dbg_adr = 32'h225e8; force soc.dbg_do = 32'h00030713; #1000;
force soc.dbg_adr = 32'h225ec; force soc.dbg_do = 32'h070e0513; #1000;
force soc.dbg_adr = 32'h225f0; force soc.dbg_do = 32'h00112e23; #1000;
force soc.dbg_adr = 32'h225f4; force soc.dbg_do = 32'h02f12a23; #1000;
force soc.dbg_adr = 32'h225f8; force soc.dbg_do = 32'h03012c23; #1000;
force soc.dbg_adr = 32'h225fc; force soc.dbg_do = 32'h03112e23; #1000;
force soc.dbg_adr = 32'h22600; force soc.dbg_do = 32'h00612623; #1000;
force soc.dbg_adr = 32'h22604; force soc.dbg_do = 32'hfd9fe0ef; #1000;
force soc.dbg_adr = 32'h22608; force soc.dbg_do = 32'h01c12083; #1000;
force soc.dbg_adr = 32'h2260c; force soc.dbg_do = 32'h04010113; #1000;
force soc.dbg_adr = 32'h22610; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h22614; force soc.dbg_do = 32'hfe010113; #1000;
force soc.dbg_adr = 32'h22618; force soc.dbg_do = 32'h00050693; #1000;
force soc.dbg_adr = 32'h2261c; force soc.dbg_do = 32'h00021537; #1000;
force soc.dbg_adr = 32'h22620; force soc.dbg_do = 32'h00058713; #1000;
force soc.dbg_adr = 32'h22624; force soc.dbg_do = 32'h5bc50513; #1000;
force soc.dbg_adr = 32'h22628; force soc.dbg_do = 32'h00c10593; #1000;
force soc.dbg_adr = 32'h2262c; force soc.dbg_do = 32'hfff00613; #1000;
force soc.dbg_adr = 32'h22630; force soc.dbg_do = 32'h00112e23; #1000;
force soc.dbg_adr = 32'h22634; force soc.dbg_do = 32'hfa9fe0ef; #1000;
force soc.dbg_adr = 32'h22638; force soc.dbg_do = 32'h01c12083; #1000;
force soc.dbg_adr = 32'h2263c; force soc.dbg_do = 32'h02010113; #1000;
force soc.dbg_adr = 32'h22640; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h22644; force soc.dbg_do = 32'h00058893; #1000;
force soc.dbg_adr = 32'h22648; force soc.dbg_do = 32'h00060813; #1000;
force soc.dbg_adr = 32'h2264c; force soc.dbg_do = 32'h000217b7; #1000;
force soc.dbg_adr = 32'h22650; force soc.dbg_do = 32'h00068713; #1000;
force soc.dbg_adr = 32'h22654; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h22658; force soc.dbg_do = 32'h00088613; #1000;
force soc.dbg_adr = 32'h2265c; force soc.dbg_do = 32'h00080693; #1000;
force soc.dbg_adr = 32'h22660; force soc.dbg_do = 32'h07078513; #1000;
force soc.dbg_adr = 32'h22664; force soc.dbg_do = 32'hf79fe06f; #1000;
force soc.dbg_adr = 32'h22668; force soc.dbg_do = 32'hfc010113; #1000;
force soc.dbg_adr = 32'h2266c; force soc.dbg_do = 32'h02c10313; #1000;
force soc.dbg_adr = 32'h22670; force soc.dbg_do = 32'h00021f37; #1000;
force soc.dbg_adr = 32'h22674; force soc.dbg_do = 32'h00050e93; #1000;
force soc.dbg_adr = 32'h22678; force soc.dbg_do = 32'h00058e13; #1000;
force soc.dbg_adr = 32'h2267c; force soc.dbg_do = 32'h02d12623; #1000;
force soc.dbg_adr = 32'h22680; force soc.dbg_do = 32'h02e12823; #1000;
force soc.dbg_adr = 32'h22684; force soc.dbg_do = 32'h00060693; #1000;
force soc.dbg_adr = 32'h22688; force soc.dbg_do = 32'h00810593; #1000;
force soc.dbg_adr = 32'h2268c; force soc.dbg_do = 32'h00030713; #1000;
force soc.dbg_adr = 32'h22690; force soc.dbg_do = 32'h5c8f0513; #1000;
force soc.dbg_adr = 32'h22694; force soc.dbg_do = 32'hfff00613; #1000;
force soc.dbg_adr = 32'h22698; force soc.dbg_do = 32'h00112e23; #1000;
force soc.dbg_adr = 32'h2269c; force soc.dbg_do = 32'h01d12423; #1000;
force soc.dbg_adr = 32'h226a0; force soc.dbg_do = 32'h01c12623; #1000;
force soc.dbg_adr = 32'h226a4; force soc.dbg_do = 32'h02f12a23; #1000;
force soc.dbg_adr = 32'h226a8; force soc.dbg_do = 32'h03012c23; #1000;
force soc.dbg_adr = 32'h226ac; force soc.dbg_do = 32'h03112e23; #1000;
force soc.dbg_adr = 32'h226b0; force soc.dbg_do = 32'h00612223; #1000;
force soc.dbg_adr = 32'h226b4; force soc.dbg_do = 32'hf29fe0ef; #1000;
force soc.dbg_adr = 32'h226b8; force soc.dbg_do = 32'h01c12083; #1000;
force soc.dbg_adr = 32'h226bc; force soc.dbg_do = 32'h04010113; #1000;
force soc.dbg_adr = 32'h226c0; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h226c4; force soc.dbg_do = 32'hfd010113; #1000;
force soc.dbg_adr = 32'h226c8; force soc.dbg_do = 32'h01412c23; #1000;
force soc.dbg_adr = 32'h226cc; force soc.dbg_do = 32'h02112623; #1000;
force soc.dbg_adr = 32'h226d0; force soc.dbg_do = 32'h02812423; #1000;
force soc.dbg_adr = 32'h226d4; force soc.dbg_do = 32'h02912223; #1000;
force soc.dbg_adr = 32'h226d8; force soc.dbg_do = 32'h03212023; #1000;
force soc.dbg_adr = 32'h226dc; force soc.dbg_do = 32'h01312e23; #1000;
force soc.dbg_adr = 32'h226e0; force soc.dbg_do = 32'h01512a23; #1000;
force soc.dbg_adr = 32'h226e4; force soc.dbg_do = 32'h01612823; #1000;
force soc.dbg_adr = 32'h226e8; force soc.dbg_do = 32'h01712623; #1000;
force soc.dbg_adr = 32'h226ec; force soc.dbg_do = 32'h01812423; #1000;
force soc.dbg_adr = 32'h226f0; force soc.dbg_do = 32'h01912223; #1000;
force soc.dbg_adr = 32'h226f4; force soc.dbg_do = 32'h01a12023; #1000;
force soc.dbg_adr = 32'h226f8; force soc.dbg_do = 32'h00050a13; #1000;
force soc.dbg_adr = 32'h226fc; force soc.dbg_do = 32'h38069663; #1000;
force soc.dbg_adr = 32'h22700; force soc.dbg_do = 32'h000247b7; #1000;
force soc.dbg_adr = 32'h22704; force soc.dbg_do = 32'h00060993; #1000;
force soc.dbg_adr = 32'h22708; force soc.dbg_do = 32'h00050493; #1000;
force soc.dbg_adr = 32'h2270c; force soc.dbg_do = 32'h20878793; #1000;
force soc.dbg_adr = 32'h22710; force soc.dbg_do = 32'h12c5f863; #1000;
force soc.dbg_adr = 32'h22714; force soc.dbg_do = 32'h00010737; #1000;
force soc.dbg_adr = 32'h22718; force soc.dbg_do = 32'h00058913; #1000;
force soc.dbg_adr = 32'h2271c; force soc.dbg_do = 32'h10e67863; #1000;
force soc.dbg_adr = 32'h22720; force soc.dbg_do = 32'h10063713; #1000;
force soc.dbg_adr = 32'h22724; force soc.dbg_do = 32'h00173713; #1000;
force soc.dbg_adr = 32'h22728; force soc.dbg_do = 32'h00371713; #1000;
force soc.dbg_adr = 32'h2272c; force soc.dbg_do = 32'h00e656b3; #1000;
force soc.dbg_adr = 32'h22730; force soc.dbg_do = 32'h00d787b3; #1000;
force soc.dbg_adr = 32'h22734; force soc.dbg_do = 32'h0007c783; #1000;
force soc.dbg_adr = 32'h22738; force soc.dbg_do = 32'h02000693; #1000;
force soc.dbg_adr = 32'h2273c; force soc.dbg_do = 32'h00e787b3; #1000;
force soc.dbg_adr = 32'h22740; force soc.dbg_do = 32'h40f68733; #1000;
force soc.dbg_adr = 32'h22744; force soc.dbg_do = 32'h00f68c63; #1000;
force soc.dbg_adr = 32'h22748; force soc.dbg_do = 32'h00e59933; #1000;
force soc.dbg_adr = 32'h2274c; force soc.dbg_do = 32'h00fa57b3; #1000;
force soc.dbg_adr = 32'h22750; force soc.dbg_do = 32'h00e619b3; #1000;
force soc.dbg_adr = 32'h22754; force soc.dbg_do = 32'h0127e933; #1000;
force soc.dbg_adr = 32'h22758; force soc.dbg_do = 32'h00ea14b3; #1000;
force soc.dbg_adr = 32'h2275c; force soc.dbg_do = 32'h0109da93; #1000;
force soc.dbg_adr = 32'h22760; force soc.dbg_do = 32'h000a8593; #1000;
force soc.dbg_adr = 32'h22764; force soc.dbg_do = 32'h00090513; #1000;
force soc.dbg_adr = 32'h22768; force soc.dbg_do = 32'h01099b13; #1000;
force soc.dbg_adr = 32'h2276c; force soc.dbg_do = 32'h310010ef; #1000;
force soc.dbg_adr = 32'h22770; force soc.dbg_do = 32'h010b5b13; #1000;
force soc.dbg_adr = 32'h22774; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h22778; force soc.dbg_do = 32'h00050a13; #1000;
force soc.dbg_adr = 32'h2277c; force soc.dbg_do = 32'h000b0513; #1000;
force soc.dbg_adr = 32'h22780; force soc.dbg_do = 32'h2d0010ef; #1000;
force soc.dbg_adr = 32'h22784; force soc.dbg_do = 32'h00050413; #1000;
force soc.dbg_adr = 32'h22788; force soc.dbg_do = 32'h000a8593; #1000;
force soc.dbg_adr = 32'h2278c; force soc.dbg_do = 32'h00090513; #1000;
force soc.dbg_adr = 32'h22790; force soc.dbg_do = 32'h334010ef; #1000;
force soc.dbg_adr = 32'h22794; force soc.dbg_do = 32'h01051513; #1000;
force soc.dbg_adr = 32'h22798; force soc.dbg_do = 32'h0104d713; #1000;
force soc.dbg_adr = 32'h2279c; force soc.dbg_do = 32'h00a76733; #1000;
force soc.dbg_adr = 32'h227a0; force soc.dbg_do = 32'h000a0913; #1000;
force soc.dbg_adr = 32'h227a4; force soc.dbg_do = 32'h00877e63; #1000;
force soc.dbg_adr = 32'h227a8; force soc.dbg_do = 32'h00e98733; #1000;
force soc.dbg_adr = 32'h227ac; force soc.dbg_do = 32'hfffa0913; #1000;
force soc.dbg_adr = 32'h227b0; force soc.dbg_do = 32'h01376863; #1000;
force soc.dbg_adr = 32'h227b4; force soc.dbg_do = 32'h00877663; #1000;
force soc.dbg_adr = 32'h227b8; force soc.dbg_do = 32'hffea0913; #1000;
force soc.dbg_adr = 32'h227bc; force soc.dbg_do = 32'h01370733; #1000;
force soc.dbg_adr = 32'h227c0; force soc.dbg_do = 32'h40870433; #1000;
force soc.dbg_adr = 32'h227c4; force soc.dbg_do = 32'h000a8593; #1000;
force soc.dbg_adr = 32'h227c8; force soc.dbg_do = 32'h00040513; #1000;
force soc.dbg_adr = 32'h227cc; force soc.dbg_do = 32'h2b0010ef; #1000;
force soc.dbg_adr = 32'h227d0; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h227d4; force soc.dbg_do = 32'h00050a13; #1000;
force soc.dbg_adr = 32'h227d8; force soc.dbg_do = 32'h000b0513; #1000;
force soc.dbg_adr = 32'h227dc; force soc.dbg_do = 32'h274010ef; #1000;
force soc.dbg_adr = 32'h227e0; force soc.dbg_do = 32'h00050b13; #1000;
force soc.dbg_adr = 32'h227e4; force soc.dbg_do = 32'h000a8593; #1000;
force soc.dbg_adr = 32'h227e8; force soc.dbg_do = 32'h00040513; #1000;
force soc.dbg_adr = 32'h227ec; force soc.dbg_do = 32'h2d8010ef; #1000;
force soc.dbg_adr = 32'h227f0; force soc.dbg_do = 32'h01049493; #1000;
force soc.dbg_adr = 32'h227f4; force soc.dbg_do = 32'h01051513; #1000;
force soc.dbg_adr = 32'h227f8; force soc.dbg_do = 32'h0104d493; #1000;
force soc.dbg_adr = 32'h227fc; force soc.dbg_do = 32'h00a4e4b3; #1000;
force soc.dbg_adr = 32'h22800; force soc.dbg_do = 32'h000a0713; #1000;
force soc.dbg_adr = 32'h22804; force soc.dbg_do = 32'h0164fc63; #1000;
force soc.dbg_adr = 32'h22808; force soc.dbg_do = 32'h009984b3; #1000;
force soc.dbg_adr = 32'h2280c; force soc.dbg_do = 32'hfffa0713; #1000;
force soc.dbg_adr = 32'h22810; force soc.dbg_do = 32'h0134e663; #1000;
force soc.dbg_adr = 32'h22814; force soc.dbg_do = 32'h0164f463; #1000;
force soc.dbg_adr = 32'h22818; force soc.dbg_do = 32'hffea0713; #1000;
force soc.dbg_adr = 32'h2281c; force soc.dbg_do = 32'h01091793; #1000;
force soc.dbg_adr = 32'h22820; force soc.dbg_do = 32'h00e7e7b3; #1000;
force soc.dbg_adr = 32'h22824; force soc.dbg_do = 32'h00000913; #1000;
force soc.dbg_adr = 32'h22828; force soc.dbg_do = 32'h1200006f; #1000;
force soc.dbg_adr = 32'h2282c; force soc.dbg_do = 32'h010006b7; #1000;
force soc.dbg_adr = 32'h22830; force soc.dbg_do = 32'h01800713; #1000;
force soc.dbg_adr = 32'h22834; force soc.dbg_do = 32'heed67ce3; #1000;
force soc.dbg_adr = 32'h22838; force soc.dbg_do = 32'h01000713; #1000;
force soc.dbg_adr = 32'h2283c; force soc.dbg_do = 32'hef1ff06f; #1000;
force soc.dbg_adr = 32'h22840; force soc.dbg_do = 32'h00000713; #1000;
force soc.dbg_adr = 32'h22844; force soc.dbg_do = 32'h00060c63; #1000;
force soc.dbg_adr = 32'h22848; force soc.dbg_do = 32'h00010737; #1000;
force soc.dbg_adr = 32'h2284c; force soc.dbg_do = 32'h12e67e63; #1000;
force soc.dbg_adr = 32'h22850; force soc.dbg_do = 32'h10063713; #1000;
force soc.dbg_adr = 32'h22854; force soc.dbg_do = 32'h00173713; #1000;
force soc.dbg_adr = 32'h22858; force soc.dbg_do = 32'h00371713; #1000;
force soc.dbg_adr = 32'h2285c; force soc.dbg_do = 32'h00e656b3; #1000;
force soc.dbg_adr = 32'h22860; force soc.dbg_do = 32'h00d787b3; #1000;
force soc.dbg_adr = 32'h22864; force soc.dbg_do = 32'h0007c783; #1000;
force soc.dbg_adr = 32'h22868; force soc.dbg_do = 32'h02000693; #1000;
force soc.dbg_adr = 32'h2286c; force soc.dbg_do = 32'h00e787b3; #1000;
force soc.dbg_adr = 32'h22870; force soc.dbg_do = 32'h40f68733; #1000;
force soc.dbg_adr = 32'h22874; force soc.dbg_do = 32'h12f69463; #1000;
force soc.dbg_adr = 32'h22878; force soc.dbg_do = 32'h40c58a33; #1000;
force soc.dbg_adr = 32'h2287c; force soc.dbg_do = 32'h00100913; #1000;
force soc.dbg_adr = 32'h22880; force soc.dbg_do = 32'h0109db13; #1000;
force soc.dbg_adr = 32'h22884; force soc.dbg_do = 32'h000b0593; #1000;
force soc.dbg_adr = 32'h22888; force soc.dbg_do = 32'h000a0513; #1000;
force soc.dbg_adr = 32'h2288c; force soc.dbg_do = 32'h01099b93; #1000;
force soc.dbg_adr = 32'h22890; force soc.dbg_do = 32'h1ec010ef; #1000;
force soc.dbg_adr = 32'h22894; force soc.dbg_do = 32'h010bdb93; #1000;
force soc.dbg_adr = 32'h22898; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h2289c; force soc.dbg_do = 32'h00050c13; #1000;
force soc.dbg_adr = 32'h228a0; force soc.dbg_do = 32'h000b8513; #1000;
force soc.dbg_adr = 32'h228a4; force soc.dbg_do = 32'h1ac010ef; #1000;
force soc.dbg_adr = 32'h228a8; force soc.dbg_do = 32'h00050a93; #1000;
force soc.dbg_adr = 32'h228ac; force soc.dbg_do = 32'h000b0593; #1000;
force soc.dbg_adr = 32'h228b0; force soc.dbg_do = 32'h000a0513; #1000;
force soc.dbg_adr = 32'h228b4; force soc.dbg_do = 32'h210010ef; #1000;
force soc.dbg_adr = 32'h228b8; force soc.dbg_do = 32'h01051513; #1000;
force soc.dbg_adr = 32'h228bc; force soc.dbg_do = 32'h0104d713; #1000;
force soc.dbg_adr = 32'h228c0; force soc.dbg_do = 32'h00a76733; #1000;
force soc.dbg_adr = 32'h228c4; force soc.dbg_do = 32'h000c0a13; #1000;
force soc.dbg_adr = 32'h228c8; force soc.dbg_do = 32'h01577e63; #1000;
force soc.dbg_adr = 32'h228cc; force soc.dbg_do = 32'h00e98733; #1000;
force soc.dbg_adr = 32'h228d0; force soc.dbg_do = 32'hfffc0a13; #1000;
force soc.dbg_adr = 32'h228d4; force soc.dbg_do = 32'h01376863; #1000;
force soc.dbg_adr = 32'h228d8; force soc.dbg_do = 32'h01577663; #1000;
force soc.dbg_adr = 32'h228dc; force soc.dbg_do = 32'hffec0a13; #1000;
force soc.dbg_adr = 32'h228e0; force soc.dbg_do = 32'h01370733; #1000;
force soc.dbg_adr = 32'h228e4; force soc.dbg_do = 32'h41570433; #1000;
force soc.dbg_adr = 32'h228e8; force soc.dbg_do = 32'h000b0593; #1000;
force soc.dbg_adr = 32'h228ec; force soc.dbg_do = 32'h00040513; #1000;
force soc.dbg_adr = 32'h228f0; force soc.dbg_do = 32'h18c010ef; #1000;
force soc.dbg_adr = 32'h228f4; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h228f8; force soc.dbg_do = 32'h00050a93; #1000;
force soc.dbg_adr = 32'h228fc; force soc.dbg_do = 32'h000b8513; #1000;
force soc.dbg_adr = 32'h22900; force soc.dbg_do = 32'h150010ef; #1000;
force soc.dbg_adr = 32'h22904; force soc.dbg_do = 32'h00050b93; #1000;
force soc.dbg_adr = 32'h22908; force soc.dbg_do = 32'h000b0593; #1000;
force soc.dbg_adr = 32'h2290c; force soc.dbg_do = 32'h00040513; #1000;
force soc.dbg_adr = 32'h22910; force soc.dbg_do = 32'h1b4010ef; #1000;
force soc.dbg_adr = 32'h22914; force soc.dbg_do = 32'h01049493; #1000;
force soc.dbg_adr = 32'h22918; force soc.dbg_do = 32'h01051513; #1000;
force soc.dbg_adr = 32'h2291c; force soc.dbg_do = 32'h0104d493; #1000;
force soc.dbg_adr = 32'h22920; force soc.dbg_do = 32'h00a4e4b3; #1000;
force soc.dbg_adr = 32'h22924; force soc.dbg_do = 32'h000a8713; #1000;
force soc.dbg_adr = 32'h22928; force soc.dbg_do = 32'h0174fc63; #1000;
force soc.dbg_adr = 32'h2292c; force soc.dbg_do = 32'h009984b3; #1000;
force soc.dbg_adr = 32'h22930; force soc.dbg_do = 32'hfffa8713; #1000;
force soc.dbg_adr = 32'h22934; force soc.dbg_do = 32'h0134e663; #1000;
force soc.dbg_adr = 32'h22938; force soc.dbg_do = 32'h0174f463; #1000;
force soc.dbg_adr = 32'h2293c; force soc.dbg_do = 32'hffea8713; #1000;
force soc.dbg_adr = 32'h22940; force soc.dbg_do = 32'h010a1793; #1000;
force soc.dbg_adr = 32'h22944; force soc.dbg_do = 32'h00e7e7b3; #1000;
force soc.dbg_adr = 32'h22948; force soc.dbg_do = 32'h02c12083; #1000;
force soc.dbg_adr = 32'h2294c; force soc.dbg_do = 32'h02812403; #1000;
force soc.dbg_adr = 32'h22950; force soc.dbg_do = 32'h02412483; #1000;
force soc.dbg_adr = 32'h22954; force soc.dbg_do = 32'h01c12983; #1000;
force soc.dbg_adr = 32'h22958; force soc.dbg_do = 32'h01812a03; #1000;
force soc.dbg_adr = 32'h2295c; force soc.dbg_do = 32'h01412a83; #1000;
force soc.dbg_adr = 32'h22960; force soc.dbg_do = 32'h01012b03; #1000;
force soc.dbg_adr = 32'h22964; force soc.dbg_do = 32'h00c12b83; #1000;
force soc.dbg_adr = 32'h22968; force soc.dbg_do = 32'h00812c03; #1000;
force soc.dbg_adr = 32'h2296c; force soc.dbg_do = 32'h00412c83; #1000;
force soc.dbg_adr = 32'h22970; force soc.dbg_do = 32'h00012d03; #1000;
force soc.dbg_adr = 32'h22974; force soc.dbg_do = 32'h00090593; #1000;
force soc.dbg_adr = 32'h22978; force soc.dbg_do = 32'h00078513; #1000;
force soc.dbg_adr = 32'h2297c; force soc.dbg_do = 32'h02012903; #1000;
force soc.dbg_adr = 32'h22980; force soc.dbg_do = 32'h03010113; #1000;
force soc.dbg_adr = 32'h22984; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h22988; force soc.dbg_do = 32'h010006b7; #1000;
force soc.dbg_adr = 32'h2298c; force soc.dbg_do = 32'h01800713; #1000;
force soc.dbg_adr = 32'h22990; force soc.dbg_do = 32'hecd676e3; #1000;
force soc.dbg_adr = 32'h22994; force soc.dbg_do = 32'h01000713; #1000;
force soc.dbg_adr = 32'h22998; force soc.dbg_do = 32'hec5ff06f; #1000;
force soc.dbg_adr = 32'h2299c; force soc.dbg_do = 32'h00e619b3; #1000;
force soc.dbg_adr = 32'h229a0; force soc.dbg_do = 32'h00f5d933; #1000;
force soc.dbg_adr = 32'h229a4; force soc.dbg_do = 32'h0109db93; #1000;
force soc.dbg_adr = 32'h229a8; force soc.dbg_do = 32'h00e595b3; #1000;
force soc.dbg_adr = 32'h229ac; force soc.dbg_do = 32'h00fa57b3; #1000;
force soc.dbg_adr = 32'h229b0; force soc.dbg_do = 32'h00b7eab3; #1000;
force soc.dbg_adr = 32'h229b4; force soc.dbg_do = 32'h00ea14b3; #1000;
force soc.dbg_adr = 32'h229b8; force soc.dbg_do = 32'h000b8593; #1000;
force soc.dbg_adr = 32'h229bc; force soc.dbg_do = 32'h00090513; #1000;
force soc.dbg_adr = 32'h229c0; force soc.dbg_do = 32'h01099a13; #1000;
force soc.dbg_adr = 32'h229c4; force soc.dbg_do = 32'h0b8010ef; #1000;
force soc.dbg_adr = 32'h229c8; force soc.dbg_do = 32'h010a5a13; #1000;
force soc.dbg_adr = 32'h229cc; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h229d0; force soc.dbg_do = 32'h00050b13; #1000;
force soc.dbg_adr = 32'h229d4; force soc.dbg_do = 32'h000a0513; #1000;
force soc.dbg_adr = 32'h229d8; force soc.dbg_do = 32'h078010ef; #1000;
force soc.dbg_adr = 32'h229dc; force soc.dbg_do = 32'h00050413; #1000;
force soc.dbg_adr = 32'h229e0; force soc.dbg_do = 32'h000b8593; #1000;
force soc.dbg_adr = 32'h229e4; force soc.dbg_do = 32'h00090513; #1000;
force soc.dbg_adr = 32'h229e8; force soc.dbg_do = 32'h0dc010ef; #1000;
force soc.dbg_adr = 32'h229ec; force soc.dbg_do = 32'h01051513; #1000;
force soc.dbg_adr = 32'h229f0; force soc.dbg_do = 32'h010ad713; #1000;
force soc.dbg_adr = 32'h229f4; force soc.dbg_do = 32'h00a76733; #1000;
force soc.dbg_adr = 32'h229f8; force soc.dbg_do = 32'h000b0913; #1000;
force soc.dbg_adr = 32'h229fc; force soc.dbg_do = 32'h00877e63; #1000;
force soc.dbg_adr = 32'h22a00; force soc.dbg_do = 32'h00e98733; #1000;
force soc.dbg_adr = 32'h22a04; force soc.dbg_do = 32'hfffb0913; #1000;
force soc.dbg_adr = 32'h22a08; force soc.dbg_do = 32'h01376863; #1000;
force soc.dbg_adr = 32'h22a0c; force soc.dbg_do = 32'h00877663; #1000;
force soc.dbg_adr = 32'h22a10; force soc.dbg_do = 32'hffeb0913; #1000;
force soc.dbg_adr = 32'h22a14; force soc.dbg_do = 32'h01370733; #1000;
force soc.dbg_adr = 32'h22a18; force soc.dbg_do = 32'h40870433; #1000;
force soc.dbg_adr = 32'h22a1c; force soc.dbg_do = 32'h000b8593; #1000;
force soc.dbg_adr = 32'h22a20; force soc.dbg_do = 32'h00040513; #1000;
force soc.dbg_adr = 32'h22a24; force soc.dbg_do = 32'h058010ef; #1000;
force soc.dbg_adr = 32'h22a28; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h22a2c; force soc.dbg_do = 32'h00050b13; #1000;
force soc.dbg_adr = 32'h22a30; force soc.dbg_do = 32'h000a0513; #1000;
force soc.dbg_adr = 32'h22a34; force soc.dbg_do = 32'h01c010ef; #1000;
force soc.dbg_adr = 32'h22a38; force soc.dbg_do = 32'h00050a13; #1000;
force soc.dbg_adr = 32'h22a3c; force soc.dbg_do = 32'h000b8593; #1000;
force soc.dbg_adr = 32'h22a40; force soc.dbg_do = 32'h00040513; #1000;
force soc.dbg_adr = 32'h22a44; force soc.dbg_do = 32'h080010ef; #1000;
force soc.dbg_adr = 32'h22a48; force soc.dbg_do = 32'h010a9793; #1000;
force soc.dbg_adr = 32'h22a4c; force soc.dbg_do = 32'h01051513; #1000;
force soc.dbg_adr = 32'h22a50; force soc.dbg_do = 32'h0107d793; #1000;
force soc.dbg_adr = 32'h22a54; force soc.dbg_do = 32'h00a7e7b3; #1000;
force soc.dbg_adr = 32'h22a58; force soc.dbg_do = 32'h000b0713; #1000;
force soc.dbg_adr = 32'h22a5c; force soc.dbg_do = 32'h0147fe63; #1000;
force soc.dbg_adr = 32'h22a60; force soc.dbg_do = 32'h00f987b3; #1000;
force soc.dbg_adr = 32'h22a64; force soc.dbg_do = 32'hfffb0713; #1000;
force soc.dbg_adr = 32'h22a68; force soc.dbg_do = 32'h0137e863; #1000;
force soc.dbg_adr = 32'h22a6c; force soc.dbg_do = 32'h0147f663; #1000;
force soc.dbg_adr = 32'h22a70; force soc.dbg_do = 32'hffeb0713; #1000;
force soc.dbg_adr = 32'h22a74; force soc.dbg_do = 32'h013787b3; #1000;
force soc.dbg_adr = 32'h22a78; force soc.dbg_do = 32'h01091913; #1000;
force soc.dbg_adr = 32'h22a7c; force soc.dbg_do = 32'h41478a33; #1000;
force soc.dbg_adr = 32'h22a80; force soc.dbg_do = 32'h00e96933; #1000;
force soc.dbg_adr = 32'h22a84; force soc.dbg_do = 32'hdfdff06f; #1000;
force soc.dbg_adr = 32'h22a88; force soc.dbg_do = 32'h1ed5ec63; #1000;
force soc.dbg_adr = 32'h22a8c; force soc.dbg_do = 32'h000107b7; #1000;
force soc.dbg_adr = 32'h22a90; force soc.dbg_do = 32'h04f6f463; #1000;
force soc.dbg_adr = 32'h22a94; force soc.dbg_do = 32'h1006b713; #1000;
force soc.dbg_adr = 32'h22a98; force soc.dbg_do = 32'h00173713; #1000;
force soc.dbg_adr = 32'h22a9c; force soc.dbg_do = 32'h00371713; #1000;
force soc.dbg_adr = 32'h22aa0; force soc.dbg_do = 32'h000247b7; #1000;
force soc.dbg_adr = 32'h22aa4; force soc.dbg_do = 32'h00e6d533; #1000;
force soc.dbg_adr = 32'h22aa8; force soc.dbg_do = 32'h20878793; #1000;
force soc.dbg_adr = 32'h22aac; force soc.dbg_do = 32'h00a787b3; #1000;
force soc.dbg_adr = 32'h22ab0; force soc.dbg_do = 32'h0007c803; #1000;
force soc.dbg_adr = 32'h22ab4; force soc.dbg_do = 32'h02000793; #1000;
force soc.dbg_adr = 32'h22ab8; force soc.dbg_do = 32'h00e80833; #1000;
force soc.dbg_adr = 32'h22abc; force soc.dbg_do = 32'h41078933; #1000;
force soc.dbg_adr = 32'h22ac0; force soc.dbg_do = 32'h03079663; #1000;
force soc.dbg_adr = 32'h22ac4; force soc.dbg_do = 32'h00100793; #1000;
force soc.dbg_adr = 32'h22ac8; force soc.dbg_do = 32'he8b6e0e3; #1000;
force soc.dbg_adr = 32'h22acc; force soc.dbg_do = 32'h00ca37b3; #1000;
force soc.dbg_adr = 32'h22ad0; force soc.dbg_do = 32'h0017b793; #1000;
force soc.dbg_adr = 32'h22ad4; force soc.dbg_do = 32'he75ff06f; #1000;
force soc.dbg_adr = 32'h22ad8; force soc.dbg_do = 32'h010007b7; #1000;
force soc.dbg_adr = 32'h22adc; force soc.dbg_do = 32'h01800713; #1000;
force soc.dbg_adr = 32'h22ae0; force soc.dbg_do = 32'hfcf6f0e3; #1000;
force soc.dbg_adr = 32'h22ae4; force soc.dbg_do = 32'h01000713; #1000;
force soc.dbg_adr = 32'h22ae8; force soc.dbg_do = 32'hfb9ff06f; #1000;
force soc.dbg_adr = 32'h22aec; force soc.dbg_do = 32'h012696b3; #1000;
force soc.dbg_adr = 32'h22af0; force soc.dbg_do = 32'h01065ab3; #1000;
force soc.dbg_adr = 32'h22af4; force soc.dbg_do = 32'h00daeab3; #1000;
force soc.dbg_adr = 32'h22af8; force soc.dbg_do = 32'h0105d9b3; #1000;
force soc.dbg_adr = 32'h22afc; force soc.dbg_do = 32'h010adc13; #1000;
force soc.dbg_adr = 32'h22b00; force soc.dbg_do = 32'h010a5833; #1000;
force soc.dbg_adr = 32'h22b04; force soc.dbg_do = 32'h012595b3; #1000;
force soc.dbg_adr = 32'h22b08; force soc.dbg_do = 32'h00b864b3; #1000;
force soc.dbg_adr = 32'h22b0c; force soc.dbg_do = 32'h010a9b93; #1000;
force soc.dbg_adr = 32'h22b10; force soc.dbg_do = 32'h000c0593; #1000;
force soc.dbg_adr = 32'h22b14; force soc.dbg_do = 32'h00098513; #1000;
force soc.dbg_adr = 32'h22b18; force soc.dbg_do = 32'h01261433; #1000;
force soc.dbg_adr = 32'h22b1c; force soc.dbg_do = 32'h010bdb93; #1000;
force soc.dbg_adr = 32'h22b20; force soc.dbg_do = 32'h75d000ef; #1000;
force soc.dbg_adr = 32'h22b24; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h22b28; force soc.dbg_do = 32'h00050d13; #1000;
force soc.dbg_adr = 32'h22b2c; force soc.dbg_do = 32'h000b8513; #1000;
force soc.dbg_adr = 32'h22b30; force soc.dbg_do = 32'h721000ef; #1000;
force soc.dbg_adr = 32'h22b34; force soc.dbg_do = 32'h00050c93; #1000;
force soc.dbg_adr = 32'h22b38; force soc.dbg_do = 32'h000c0593; #1000;
force soc.dbg_adr = 32'h22b3c; force soc.dbg_do = 32'h00098513; #1000;
force soc.dbg_adr = 32'h22b40; force soc.dbg_do = 32'h785000ef; #1000;
force soc.dbg_adr = 32'h22b44; force soc.dbg_do = 32'h01051513; #1000;
force soc.dbg_adr = 32'h22b48; force soc.dbg_do = 32'h0104d693; #1000;
force soc.dbg_adr = 32'h22b4c; force soc.dbg_do = 32'h00a6e6b3; #1000;
force soc.dbg_adr = 32'h22b50; force soc.dbg_do = 32'h000d0b13; #1000;
force soc.dbg_adr = 32'h22b54; force soc.dbg_do = 32'h0196fe63; #1000;
force soc.dbg_adr = 32'h22b58; force soc.dbg_do = 32'h00da86b3; #1000;
force soc.dbg_adr = 32'h22b5c; force soc.dbg_do = 32'hfffd0b13; #1000;
force soc.dbg_adr = 32'h22b60; force soc.dbg_do = 32'h0156e863; #1000;
force soc.dbg_adr = 32'h22b64; force soc.dbg_do = 32'h0196f663; #1000;
force soc.dbg_adr = 32'h22b68; force soc.dbg_do = 32'hffed0b13; #1000;
force soc.dbg_adr = 32'h22b6c; force soc.dbg_do = 32'h015686b3; #1000;
force soc.dbg_adr = 32'h22b70; force soc.dbg_do = 32'h419689b3; #1000;
force soc.dbg_adr = 32'h22b74; force soc.dbg_do = 32'h000c0593; #1000;
force soc.dbg_adr = 32'h22b78; force soc.dbg_do = 32'h00098513; #1000;
force soc.dbg_adr = 32'h22b7c; force soc.dbg_do = 32'h701000ef; #1000;
force soc.dbg_adr = 32'h22b80; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h22b84; force soc.dbg_do = 32'h00050c93; #1000;
force soc.dbg_adr = 32'h22b88; force soc.dbg_do = 32'h000b8513; #1000;
force soc.dbg_adr = 32'h22b8c; force soc.dbg_do = 32'h6c5000ef; #1000;
force soc.dbg_adr = 32'h22b90; force soc.dbg_do = 32'h00050b93; #1000;
force soc.dbg_adr = 32'h22b94; force soc.dbg_do = 32'h000c0593; #1000;
force soc.dbg_adr = 32'h22b98; force soc.dbg_do = 32'h00098513; #1000;
force soc.dbg_adr = 32'h22b9c; force soc.dbg_do = 32'h729000ef; #1000;
force soc.dbg_adr = 32'h22ba0; force soc.dbg_do = 32'h01049713; #1000;
force soc.dbg_adr = 32'h22ba4; force soc.dbg_do = 32'h01051513; #1000;
force soc.dbg_adr = 32'h22ba8; force soc.dbg_do = 32'h01075713; #1000;
force soc.dbg_adr = 32'h22bac; force soc.dbg_do = 32'h00a76733; #1000;
force soc.dbg_adr = 32'h22bb0; force soc.dbg_do = 32'h000c8693; #1000;
force soc.dbg_adr = 32'h22bb4; force soc.dbg_do = 32'h01777e63; #1000;
force soc.dbg_adr = 32'h22bb8; force soc.dbg_do = 32'h00ea8733; #1000;
force soc.dbg_adr = 32'h22bbc; force soc.dbg_do = 32'hfffc8693; #1000;
force soc.dbg_adr = 32'h22bc0; force soc.dbg_do = 32'h01576863; #1000;
force soc.dbg_adr = 32'h22bc4; force soc.dbg_do = 32'h01777663; #1000;
force soc.dbg_adr = 32'h22bc8; force soc.dbg_do = 32'hffec8693; #1000;
force soc.dbg_adr = 32'h22bcc; force soc.dbg_do = 32'h01570733; #1000;
force soc.dbg_adr = 32'h22bd0; force soc.dbg_do = 32'h010b1793; #1000;
force soc.dbg_adr = 32'h22bd4; force soc.dbg_do = 32'h01069813; #1000;
force soc.dbg_adr = 32'h22bd8; force soc.dbg_do = 32'h01041313; #1000;
force soc.dbg_adr = 32'h22bdc; force soc.dbg_do = 32'h00d7e7b3; #1000;
force soc.dbg_adr = 32'h22be0; force soc.dbg_do = 32'h01085813; #1000;
force soc.dbg_adr = 32'h22be4; force soc.dbg_do = 32'h01035313; #1000;
force soc.dbg_adr = 32'h22be8; force soc.dbg_do = 32'h41770733; #1000;
force soc.dbg_adr = 32'h22bec; force soc.dbg_do = 32'h0107de13; #1000;
force soc.dbg_adr = 32'h22bf0; force soc.dbg_do = 32'h01045413; #1000;
force soc.dbg_adr = 32'h22bf4; force soc.dbg_do = 32'h00080513; #1000;
force soc.dbg_adr = 32'h22bf8; force soc.dbg_do = 32'h00030593; #1000;
force soc.dbg_adr = 32'h22bfc; force soc.dbg_do = 32'h655000ef; #1000;
force soc.dbg_adr = 32'h22c00; force soc.dbg_do = 32'h00050893; #1000;
force soc.dbg_adr = 32'h22c04; force soc.dbg_do = 32'h00040593; #1000;
force soc.dbg_adr = 32'h22c08; force soc.dbg_do = 32'h00080513; #1000;
force soc.dbg_adr = 32'h22c0c; force soc.dbg_do = 32'h645000ef; #1000;
force soc.dbg_adr = 32'h22c10; force soc.dbg_do = 32'h00050813; #1000;
force soc.dbg_adr = 32'h22c14; force soc.dbg_do = 32'h00030593; #1000;
force soc.dbg_adr = 32'h22c18; force soc.dbg_do = 32'h000e0513; #1000;
force soc.dbg_adr = 32'h22c1c; force soc.dbg_do = 32'h635000ef; #1000;
force soc.dbg_adr = 32'h22c20; force soc.dbg_do = 32'h00050313; #1000;
force soc.dbg_adr = 32'h22c24; force soc.dbg_do = 32'h00040593; #1000;
force soc.dbg_adr = 32'h22c28; force soc.dbg_do = 32'h000e0513; #1000;
force soc.dbg_adr = 32'h22c2c; force soc.dbg_do = 32'h625000ef; #1000;
force soc.dbg_adr = 32'h22c30; force soc.dbg_do = 32'h0108d693; #1000;
force soc.dbg_adr = 32'h22c34; force soc.dbg_do = 32'h00680833; #1000;
force soc.dbg_adr = 32'h22c38; force soc.dbg_do = 32'h010686b3; #1000;
force soc.dbg_adr = 32'h22c3c; force soc.dbg_do = 32'h00050613; #1000;
force soc.dbg_adr = 32'h22c40; force soc.dbg_do = 32'h0066f663; #1000;
force soc.dbg_adr = 32'h22c44; force soc.dbg_do = 32'h000105b7; #1000;
force soc.dbg_adr = 32'h22c48; force soc.dbg_do = 32'h00b50633; #1000;
force soc.dbg_adr = 32'h22c4c; force soc.dbg_do = 32'h0106d593; #1000;
force soc.dbg_adr = 32'h22c50; force soc.dbg_do = 32'h00c58633; #1000;
force soc.dbg_adr = 32'h22c54; force soc.dbg_do = 32'h02c76263; #1000;
force soc.dbg_adr = 32'h22c58; force soc.dbg_do = 32'hbcc716e3; #1000;
force soc.dbg_adr = 32'h22c5c; force soc.dbg_do = 32'h01089893; #1000;
force soc.dbg_adr = 32'h22c60; force soc.dbg_do = 32'h01069693; #1000;
force soc.dbg_adr = 32'h22c64; force soc.dbg_do = 32'h0108d893; #1000;
force soc.dbg_adr = 32'h22c68; force soc.dbg_do = 32'h012a1733; #1000;
force soc.dbg_adr = 32'h22c6c; force soc.dbg_do = 32'h011686b3; #1000;
force soc.dbg_adr = 32'h22c70; force soc.dbg_do = 32'h00000913; #1000;
force soc.dbg_adr = 32'h22c74; force soc.dbg_do = 32'hccd77ae3; #1000;
force soc.dbg_adr = 32'h22c78; force soc.dbg_do = 32'hfff78793; #1000;
force soc.dbg_adr = 32'h22c7c; force soc.dbg_do = 32'hba9ff06f; #1000;
force soc.dbg_adr = 32'h22c80; force soc.dbg_do = 32'h00000913; #1000;
force soc.dbg_adr = 32'h22c84; force soc.dbg_do = 32'h00000793; #1000;
force soc.dbg_adr = 32'h22c88; force soc.dbg_do = 32'hcc1ff06f; #1000;
force soc.dbg_adr = 32'h22c8c; force soc.dbg_do = 32'hfd010113; #1000;
force soc.dbg_adr = 32'h22c90; force soc.dbg_do = 32'h02812423; #1000;
force soc.dbg_adr = 32'h22c94; force soc.dbg_do = 32'h02912223; #1000;
force soc.dbg_adr = 32'h22c98; force soc.dbg_do = 32'h02112623; #1000;
force soc.dbg_adr = 32'h22c9c; force soc.dbg_do = 32'h03212023; #1000;
force soc.dbg_adr = 32'h22ca0; force soc.dbg_do = 32'h01312e23; #1000;
force soc.dbg_adr = 32'h22ca4; force soc.dbg_do = 32'h01412c23; #1000;
force soc.dbg_adr = 32'h22ca8; force soc.dbg_do = 32'h01512a23; #1000;
force soc.dbg_adr = 32'h22cac; force soc.dbg_do = 32'h01612823; #1000;
force soc.dbg_adr = 32'h22cb0; force soc.dbg_do = 32'h01712623; #1000;
force soc.dbg_adr = 32'h22cb4; force soc.dbg_do = 32'h01812423; #1000;
force soc.dbg_adr = 32'h22cb8; force soc.dbg_do = 32'h01912223; #1000;
force soc.dbg_adr = 32'h22cbc; force soc.dbg_do = 32'h01a12023; #1000;
force soc.dbg_adr = 32'h22cc0; force soc.dbg_do = 32'h00050413; #1000;
force soc.dbg_adr = 32'h22cc4; force soc.dbg_do = 32'h00058493; #1000;
force soc.dbg_adr = 32'h22cc8; force soc.dbg_do = 32'h24069c63; #1000;
force soc.dbg_adr = 32'h22ccc; force soc.dbg_do = 32'h000247b7; #1000;
force soc.dbg_adr = 32'h22cd0; force soc.dbg_do = 32'h00060993; #1000;
force soc.dbg_adr = 32'h22cd4; force soc.dbg_do = 32'h20878793; #1000;
force soc.dbg_adr = 32'h22cd8; force soc.dbg_do = 32'h12c5fe63; #1000;
force soc.dbg_adr = 32'h22cdc; force soc.dbg_do = 32'h00010737; #1000;
force soc.dbg_adr = 32'h22ce0; force soc.dbg_do = 32'h12e67063; #1000;
force soc.dbg_adr = 32'h22ce4; force soc.dbg_do = 32'h10063713; #1000;
force soc.dbg_adr = 32'h22ce8; force soc.dbg_do = 32'h00173713; #1000;
force soc.dbg_adr = 32'h22cec; force soc.dbg_do = 32'h00371713; #1000;
force soc.dbg_adr = 32'h22cf0; force soc.dbg_do = 32'h00e656b3; #1000;
force soc.dbg_adr = 32'h22cf4; force soc.dbg_do = 32'h00d787b3; #1000;
force soc.dbg_adr = 32'h22cf8; force soc.dbg_do = 32'h0007c783; #1000;
force soc.dbg_adr = 32'h22cfc; force soc.dbg_do = 32'h00e787b3; #1000;
force soc.dbg_adr = 32'h22d00; force soc.dbg_do = 32'h02000713; #1000;
force soc.dbg_adr = 32'h22d04; force soc.dbg_do = 32'h40f70933; #1000;
force soc.dbg_adr = 32'h22d08; force soc.dbg_do = 32'h00f70c63; #1000;
force soc.dbg_adr = 32'h22d0c; force soc.dbg_do = 32'h012594b3; #1000;
force soc.dbg_adr = 32'h22d10; force soc.dbg_do = 32'h00f557b3; #1000;
force soc.dbg_adr = 32'h22d14; force soc.dbg_do = 32'h012619b3; #1000;
force soc.dbg_adr = 32'h22d18; force soc.dbg_do = 32'h0097e4b3; #1000;
force soc.dbg_adr = 32'h22d1c; force soc.dbg_do = 32'h01251433; #1000;
force soc.dbg_adr = 32'h22d20; force soc.dbg_do = 32'h0109da93; #1000;
force soc.dbg_adr = 32'h22d24; force soc.dbg_do = 32'h000a8593; #1000;
force soc.dbg_adr = 32'h22d28; force soc.dbg_do = 32'h01099b13; #1000;
force soc.dbg_adr = 32'h22d2c; force soc.dbg_do = 32'h00048513; #1000;
force soc.dbg_adr = 32'h22d30; force soc.dbg_do = 32'h54d000ef; #1000;
force soc.dbg_adr = 32'h22d34; force soc.dbg_do = 32'h010b5b13; #1000;
force soc.dbg_adr = 32'h22d38; force soc.dbg_do = 32'h000b0593; #1000;
force soc.dbg_adr = 32'h22d3c; force soc.dbg_do = 32'h515000ef; #1000;
force soc.dbg_adr = 32'h22d40; force soc.dbg_do = 32'h00050a13; #1000;
force soc.dbg_adr = 32'h22d44; force soc.dbg_do = 32'h000a8593; #1000;
force soc.dbg_adr = 32'h22d48; force soc.dbg_do = 32'h00048513; #1000;
force soc.dbg_adr = 32'h22d4c; force soc.dbg_do = 32'h579000ef; #1000;
force soc.dbg_adr = 32'h22d50; force soc.dbg_do = 32'h01051513; #1000;
force soc.dbg_adr = 32'h22d54; force soc.dbg_do = 32'h01045793; #1000;
force soc.dbg_adr = 32'h22d58; force soc.dbg_do = 32'h00a7e7b3; #1000;
force soc.dbg_adr = 32'h22d5c; force soc.dbg_do = 32'h0147fa63; #1000;
force soc.dbg_adr = 32'h22d60; force soc.dbg_do = 32'h00f987b3; #1000;
force soc.dbg_adr = 32'h22d64; force soc.dbg_do = 32'h0137e663; #1000;
force soc.dbg_adr = 32'h22d68; force soc.dbg_do = 32'h0147f463; #1000;
force soc.dbg_adr = 32'h22d6c; force soc.dbg_do = 32'h013787b3; #1000;
force soc.dbg_adr = 32'h22d70; force soc.dbg_do = 32'h414784b3; #1000;
force soc.dbg_adr = 32'h22d74; force soc.dbg_do = 32'h000a8593; #1000;
force soc.dbg_adr = 32'h22d78; force soc.dbg_do = 32'h00048513; #1000;
force soc.dbg_adr = 32'h22d7c; force soc.dbg_do = 32'h501000ef; #1000;
force soc.dbg_adr = 32'h22d80; force soc.dbg_do = 32'h000b0593; #1000;
force soc.dbg_adr = 32'h22d84; force soc.dbg_do = 32'h4cd000ef; #1000;
force soc.dbg_adr = 32'h22d88; force soc.dbg_do = 32'h00050a13; #1000;
force soc.dbg_adr = 32'h22d8c; force soc.dbg_do = 32'h000a8593; #1000;
force soc.dbg_adr = 32'h22d90; force soc.dbg_do = 32'h00048513; #1000;
force soc.dbg_adr = 32'h22d94; force soc.dbg_do = 32'h531000ef; #1000;
force soc.dbg_adr = 32'h22d98; force soc.dbg_do = 32'h01041413; #1000;
force soc.dbg_adr = 32'h22d9c; force soc.dbg_do = 32'h01051513; #1000;
force soc.dbg_adr = 32'h22da0; force soc.dbg_do = 32'h01045413; #1000;
force soc.dbg_adr = 32'h22da4; force soc.dbg_do = 32'h00a46433; #1000;
force soc.dbg_adr = 32'h22da8; force soc.dbg_do = 32'h01447a63; #1000;
force soc.dbg_adr = 32'h22dac; force soc.dbg_do = 32'h00898433; #1000;
force soc.dbg_adr = 32'h22db0; force soc.dbg_do = 32'h01346663; #1000;
force soc.dbg_adr = 32'h22db4; force soc.dbg_do = 32'h01447463; #1000;
force soc.dbg_adr = 32'h22db8; force soc.dbg_do = 32'h01340433; #1000;
force soc.dbg_adr = 32'h22dbc; force soc.dbg_do = 32'h41440433; #1000;
force soc.dbg_adr = 32'h22dc0; force soc.dbg_do = 32'h01245533; #1000;
force soc.dbg_adr = 32'h22dc4; force soc.dbg_do = 32'h00000593; #1000;
force soc.dbg_adr = 32'h22dc8; force soc.dbg_do = 32'h02c12083; #1000;
force soc.dbg_adr = 32'h22dcc; force soc.dbg_do = 32'h02812403; #1000;
force soc.dbg_adr = 32'h22dd0; force soc.dbg_do = 32'h02412483; #1000;
force soc.dbg_adr = 32'h22dd4; force soc.dbg_do = 32'h02012903; #1000;
force soc.dbg_adr = 32'h22dd8; force soc.dbg_do = 32'h01c12983; #1000;
force soc.dbg_adr = 32'h22ddc; force soc.dbg_do = 32'h01812a03; #1000;
force soc.dbg_adr = 32'h22de0; force soc.dbg_do = 32'h01412a83; #1000;
force soc.dbg_adr = 32'h22de4; force soc.dbg_do = 32'h01012b03; #1000;
force soc.dbg_adr = 32'h22de8; force soc.dbg_do = 32'h00c12b83; #1000;
force soc.dbg_adr = 32'h22dec; force soc.dbg_do = 32'h00812c03; #1000;
force soc.dbg_adr = 32'h22df0; force soc.dbg_do = 32'h00412c83; #1000;
force soc.dbg_adr = 32'h22df4; force soc.dbg_do = 32'h00012d03; #1000;
force soc.dbg_adr = 32'h22df8; force soc.dbg_do = 32'h03010113; #1000;
force soc.dbg_adr = 32'h22dfc; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h22e00; force soc.dbg_do = 32'h010006b7; #1000;
force soc.dbg_adr = 32'h22e04; force soc.dbg_do = 32'h01800713; #1000;
force soc.dbg_adr = 32'h22e08; force soc.dbg_do = 32'heed674e3; #1000;
force soc.dbg_adr = 32'h22e0c; force soc.dbg_do = 32'h01000713; #1000;
force soc.dbg_adr = 32'h22e10; force soc.dbg_do = 32'hee1ff06f; #1000;
force soc.dbg_adr = 32'h22e14; force soc.dbg_do = 32'h00000713; #1000;
force soc.dbg_adr = 32'h22e18; force soc.dbg_do = 32'h00060c63; #1000;
force soc.dbg_adr = 32'h22e1c; force soc.dbg_do = 32'h00010737; #1000;
force soc.dbg_adr = 32'h22e20; force soc.dbg_do = 32'h0ee67663; #1000;
force soc.dbg_adr = 32'h22e24; force soc.dbg_do = 32'h10063713; #1000;
force soc.dbg_adr = 32'h22e28; force soc.dbg_do = 32'h00173713; #1000;
force soc.dbg_adr = 32'h22e2c; force soc.dbg_do = 32'h00371713; #1000;
force soc.dbg_adr = 32'h22e30; force soc.dbg_do = 32'h00e656b3; #1000;
force soc.dbg_adr = 32'h22e34; force soc.dbg_do = 32'h00d787b3; #1000;
force soc.dbg_adr = 32'h22e38; force soc.dbg_do = 32'h0007c783; #1000;
force soc.dbg_adr = 32'h22e3c; force soc.dbg_do = 32'h40c584b3; #1000;
force soc.dbg_adr = 32'h22e40; force soc.dbg_do = 32'h00e787b3; #1000;
force soc.dbg_adr = 32'h22e44; force soc.dbg_do = 32'h02000713; #1000;
force soc.dbg_adr = 32'h22e48; force soc.dbg_do = 32'h40f70933; #1000;
force soc.dbg_adr = 32'h22e4c; force soc.dbg_do = 32'hecf70ae3; #1000;
force soc.dbg_adr = 32'h22e50; force soc.dbg_do = 32'h012619b3; #1000;
force soc.dbg_adr = 32'h22e54; force soc.dbg_do = 32'h00f5dbb3; #1000;
force soc.dbg_adr = 32'h22e58; force soc.dbg_do = 32'h0109db13; #1000;
force soc.dbg_adr = 32'h22e5c; force soc.dbg_do = 32'h00f557b3; #1000;
force soc.dbg_adr = 32'h22e60; force soc.dbg_do = 32'h012595b3; #1000;
force soc.dbg_adr = 32'h22e64; force soc.dbg_do = 32'h00b7ea33; #1000;
force soc.dbg_adr = 32'h22e68; force soc.dbg_do = 32'h01251433; #1000;
force soc.dbg_adr = 32'h22e6c; force soc.dbg_do = 32'h000b0593; #1000;
force soc.dbg_adr = 32'h22e70; force soc.dbg_do = 32'h01099a93; #1000;
force soc.dbg_adr = 32'h22e74; force soc.dbg_do = 32'h000b8513; #1000;
force soc.dbg_adr = 32'h22e78; force soc.dbg_do = 32'h405000ef; #1000;
force soc.dbg_adr = 32'h22e7c; force soc.dbg_do = 32'h010ada93; #1000;
force soc.dbg_adr = 32'h22e80; force soc.dbg_do = 32'h000a8593; #1000;
force soc.dbg_adr = 32'h22e84; force soc.dbg_do = 32'h3cd000ef; #1000;
force soc.dbg_adr = 32'h22e88; force soc.dbg_do = 32'h00050493; #1000;
force soc.dbg_adr = 32'h22e8c; force soc.dbg_do = 32'h000b0593; #1000;
force soc.dbg_adr = 32'h22e90; force soc.dbg_do = 32'h000b8513; #1000;
force soc.dbg_adr = 32'h22e94; force soc.dbg_do = 32'h431000ef; #1000;
force soc.dbg_adr = 32'h22e98; force soc.dbg_do = 32'h01051513; #1000;
force soc.dbg_adr = 32'h22e9c; force soc.dbg_do = 32'h010a5713; #1000;
force soc.dbg_adr = 32'h22ea0; force soc.dbg_do = 32'h00a76733; #1000;
force soc.dbg_adr = 32'h22ea4; force soc.dbg_do = 32'h00977a63; #1000;
force soc.dbg_adr = 32'h22ea8; force soc.dbg_do = 32'h00e98733; #1000;
force soc.dbg_adr = 32'h22eac; force soc.dbg_do = 32'h01376663; #1000;
force soc.dbg_adr = 32'h22eb0; force soc.dbg_do = 32'h00977463; #1000;
force soc.dbg_adr = 32'h22eb4; force soc.dbg_do = 32'h01370733; #1000;
force soc.dbg_adr = 32'h22eb8; force soc.dbg_do = 32'h409704b3; #1000;
force soc.dbg_adr = 32'h22ebc; force soc.dbg_do = 32'h000b0593; #1000;
force soc.dbg_adr = 32'h22ec0; force soc.dbg_do = 32'h00048513; #1000;
force soc.dbg_adr = 32'h22ec4; force soc.dbg_do = 32'h3b9000ef; #1000;
force soc.dbg_adr = 32'h22ec8; force soc.dbg_do = 32'h000a8593; #1000;
force soc.dbg_adr = 32'h22ecc; force soc.dbg_do = 32'h385000ef; #1000;
force soc.dbg_adr = 32'h22ed0; force soc.dbg_do = 32'h00050a93; #1000;
force soc.dbg_adr = 32'h22ed4; force soc.dbg_do = 32'h000b0593; #1000;
force soc.dbg_adr = 32'h22ed8; force soc.dbg_do = 32'h00048513; #1000;
force soc.dbg_adr = 32'h22edc; force soc.dbg_do = 32'h3e9000ef; #1000;
force soc.dbg_adr = 32'h22ee0; force soc.dbg_do = 32'h010a1793; #1000;
force soc.dbg_adr = 32'h22ee4; force soc.dbg_do = 32'h01051513; #1000;
force soc.dbg_adr = 32'h22ee8; force soc.dbg_do = 32'h0107d793; #1000;
force soc.dbg_adr = 32'h22eec; force soc.dbg_do = 32'h00a7e7b3; #1000;
force soc.dbg_adr = 32'h22ef0; force soc.dbg_do = 32'h0157fa63; #1000;
force soc.dbg_adr = 32'h22ef4; force soc.dbg_do = 32'h00f987b3; #1000;
force soc.dbg_adr = 32'h22ef8; force soc.dbg_do = 32'h0137e663; #1000;
force soc.dbg_adr = 32'h22efc; force soc.dbg_do = 32'h0157f463; #1000;
force soc.dbg_adr = 32'h22f00; force soc.dbg_do = 32'h013787b3; #1000;
force soc.dbg_adr = 32'h22f04; force soc.dbg_do = 32'h415784b3; #1000;
force soc.dbg_adr = 32'h22f08; force soc.dbg_do = 32'he19ff06f; #1000;
force soc.dbg_adr = 32'h22f0c; force soc.dbg_do = 32'h010006b7; #1000;
force soc.dbg_adr = 32'h22f10; force soc.dbg_do = 32'h01800713; #1000;
force soc.dbg_adr = 32'h22f14; force soc.dbg_do = 32'hf0d67ee3; #1000;
force soc.dbg_adr = 32'h22f18; force soc.dbg_do = 32'h01000713; #1000;
force soc.dbg_adr = 32'h22f1c; force soc.dbg_do = 32'hf15ff06f; #1000;
force soc.dbg_adr = 32'h22f20; force soc.dbg_do = 32'head5e4e3; #1000;
force soc.dbg_adr = 32'h22f24; force soc.dbg_do = 32'h000107b7; #1000;
force soc.dbg_adr = 32'h22f28; force soc.dbg_do = 32'h04f6fe63; #1000;
force soc.dbg_adr = 32'h22f2c; force soc.dbg_do = 32'h1006b793; #1000;
force soc.dbg_adr = 32'h22f30; force soc.dbg_do = 32'h0017b793; #1000;
force soc.dbg_adr = 32'h22f34; force soc.dbg_do = 32'h00379793; #1000;
force soc.dbg_adr = 32'h22f38; force soc.dbg_do = 32'h00024737; #1000;
force soc.dbg_adr = 32'h22f3c; force soc.dbg_do = 32'h00f6d833; #1000;
force soc.dbg_adr = 32'h22f40; force soc.dbg_do = 32'h20870713; #1000;
force soc.dbg_adr = 32'h22f44; force soc.dbg_do = 32'h01070733; #1000;
force soc.dbg_adr = 32'h22f48; force soc.dbg_do = 32'h00074a83; #1000;
force soc.dbg_adr = 32'h22f4c; force soc.dbg_do = 32'h00fa8ab3; #1000;
force soc.dbg_adr = 32'h22f50; force soc.dbg_do = 32'h02000793; #1000;
force soc.dbg_adr = 32'h22f54; force soc.dbg_do = 32'h41578a33; #1000;
force soc.dbg_adr = 32'h22f58; force soc.dbg_do = 32'h05579063; #1000;
force soc.dbg_adr = 32'h22f5c; force soc.dbg_do = 32'h00b6e463; #1000;
force soc.dbg_adr = 32'h22f60; force soc.dbg_do = 32'h00c56c63; #1000;
force soc.dbg_adr = 32'h22f64; force soc.dbg_do = 32'h40c50933; #1000;
force soc.dbg_adr = 32'h22f68; force soc.dbg_do = 32'h40d586b3; #1000;
force soc.dbg_adr = 32'h22f6c; force soc.dbg_do = 32'h012534b3; #1000;
force soc.dbg_adr = 32'h22f70; force soc.dbg_do = 32'h00090413; #1000;
force soc.dbg_adr = 32'h22f74; force soc.dbg_do = 32'h409684b3; #1000;
force soc.dbg_adr = 32'h22f78; force soc.dbg_do = 32'h00040513; #1000;
force soc.dbg_adr = 32'h22f7c; force soc.dbg_do = 32'h00048593; #1000;
force soc.dbg_adr = 32'h22f80; force soc.dbg_do = 32'he49ff06f; #1000;
force soc.dbg_adr = 32'h22f84; force soc.dbg_do = 32'h01000737; #1000;
force soc.dbg_adr = 32'h22f88; force soc.dbg_do = 32'h01800793; #1000;
force soc.dbg_adr = 32'h22f8c; force soc.dbg_do = 32'hfae6f6e3; #1000;
force soc.dbg_adr = 32'h22f90; force soc.dbg_do = 32'h01000793; #1000;
force soc.dbg_adr = 32'h22f94; force soc.dbg_do = 32'hfa5ff06f; #1000;
force soc.dbg_adr = 32'h22f98; force soc.dbg_do = 32'h014696b3; #1000;
force soc.dbg_adr = 32'h22f9c; force soc.dbg_do = 32'h01565b33; #1000;
force soc.dbg_adr = 32'h22fa0; force soc.dbg_do = 32'h00db6b33; #1000;
force soc.dbg_adr = 32'h22fa4; force soc.dbg_do = 32'h0155dbb3; #1000;
force soc.dbg_adr = 32'h22fa8; force soc.dbg_do = 32'h01555433; #1000;
force soc.dbg_adr = 32'h22fac; force soc.dbg_do = 32'h014595b3; #1000;
force soc.dbg_adr = 32'h22fb0; force soc.dbg_do = 32'h010b5493; #1000;
force soc.dbg_adr = 32'h22fb4; force soc.dbg_do = 32'h00b46433; #1000;
force soc.dbg_adr = 32'h22fb8; force soc.dbg_do = 32'h014519b3; #1000;
force soc.dbg_adr = 32'h22fbc; force soc.dbg_do = 32'h00048593; #1000;
force soc.dbg_adr = 32'h22fc0; force soc.dbg_do = 32'h000b8513; #1000;
force soc.dbg_adr = 32'h22fc4; force soc.dbg_do = 32'h010b1c13; #1000;
force soc.dbg_adr = 32'h22fc8; force soc.dbg_do = 32'h01461933; #1000;
force soc.dbg_adr = 32'h22fcc; force soc.dbg_do = 32'h010c5c13; #1000;
force soc.dbg_adr = 32'h22fd0; force soc.dbg_do = 32'h2ad000ef; #1000;
force soc.dbg_adr = 32'h22fd4; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h22fd8; force soc.dbg_do = 32'h00050d13; #1000;
force soc.dbg_adr = 32'h22fdc; force soc.dbg_do = 32'h000c0513; #1000;
force soc.dbg_adr = 32'h22fe0; force soc.dbg_do = 32'h271000ef; #1000;
force soc.dbg_adr = 32'h22fe4; force soc.dbg_do = 32'h00050c93; #1000;
force soc.dbg_adr = 32'h22fe8; force soc.dbg_do = 32'h00048593; #1000;
force soc.dbg_adr = 32'h22fec; force soc.dbg_do = 32'h000b8513; #1000;
force soc.dbg_adr = 32'h22ff0; force soc.dbg_do = 32'h2d5000ef; #1000;
force soc.dbg_adr = 32'h22ff4; force soc.dbg_do = 32'h01051513; #1000;
force soc.dbg_adr = 32'h22ff8; force soc.dbg_do = 32'h01045793; #1000;
force soc.dbg_adr = 32'h22ffc; force soc.dbg_do = 32'h00a7e7b3; #1000;
force soc.dbg_adr = 32'h23000; force soc.dbg_do = 32'h000d0b93; #1000;
force soc.dbg_adr = 32'h23004; force soc.dbg_do = 32'h0197fe63; #1000;
force soc.dbg_adr = 32'h23008; force soc.dbg_do = 32'h00fb07b3; #1000;
force soc.dbg_adr = 32'h2300c; force soc.dbg_do = 32'hfffd0b93; #1000;
force soc.dbg_adr = 32'h23010; force soc.dbg_do = 32'h0167e863; #1000;
force soc.dbg_adr = 32'h23014; force soc.dbg_do = 32'h0197f663; #1000;
force soc.dbg_adr = 32'h23018; force soc.dbg_do = 32'hffed0b93; #1000;
force soc.dbg_adr = 32'h2301c; force soc.dbg_do = 32'h016787b3; #1000;
force soc.dbg_adr = 32'h23020; force soc.dbg_do = 32'h41978cb3; #1000;
force soc.dbg_adr = 32'h23024; force soc.dbg_do = 32'h00048593; #1000;
force soc.dbg_adr = 32'h23028; force soc.dbg_do = 32'h000c8513; #1000;
force soc.dbg_adr = 32'h2302c; force soc.dbg_do = 32'h251000ef; #1000;
force soc.dbg_adr = 32'h23030; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h23034; force soc.dbg_do = 32'h00050d13; #1000;
force soc.dbg_adr = 32'h23038; force soc.dbg_do = 32'h000c0513; #1000;
force soc.dbg_adr = 32'h2303c; force soc.dbg_do = 32'h215000ef; #1000;
force soc.dbg_adr = 32'h23040; force soc.dbg_do = 32'h00048593; #1000;
force soc.dbg_adr = 32'h23044; force soc.dbg_do = 32'h00050c13; #1000;
force soc.dbg_adr = 32'h23048; force soc.dbg_do = 32'h000c8513; #1000;
force soc.dbg_adr = 32'h2304c; force soc.dbg_do = 32'h279000ef; #1000;
force soc.dbg_adr = 32'h23050; force soc.dbg_do = 32'h01041593; #1000;
force soc.dbg_adr = 32'h23054; force soc.dbg_do = 32'h01051513; #1000;
force soc.dbg_adr = 32'h23058; force soc.dbg_do = 32'h0105d593; #1000;
force soc.dbg_adr = 32'h2305c; force soc.dbg_do = 32'h00a5e5b3; #1000;
force soc.dbg_adr = 32'h23060; force soc.dbg_do = 32'h000d0793; #1000;
force soc.dbg_adr = 32'h23064; force soc.dbg_do = 32'h0185fe63; #1000;
force soc.dbg_adr = 32'h23068; force soc.dbg_do = 32'h00bb05b3; #1000;
force soc.dbg_adr = 32'h2306c; force soc.dbg_do = 32'hfffd0793; #1000;
force soc.dbg_adr = 32'h23070; force soc.dbg_do = 32'h0165e863; #1000;
force soc.dbg_adr = 32'h23074; force soc.dbg_do = 32'h0185f663; #1000;
force soc.dbg_adr = 32'h23078; force soc.dbg_do = 32'hffed0793; #1000;
force soc.dbg_adr = 32'h2307c; force soc.dbg_do = 32'h016585b3; #1000;
force soc.dbg_adr = 32'h23080; force soc.dbg_do = 32'h010b9b93; #1000;
force soc.dbg_adr = 32'h23084; force soc.dbg_do = 32'h00fbebb3; #1000;
force soc.dbg_adr = 32'h23088; force soc.dbg_do = 32'h01091893; #1000;
force soc.dbg_adr = 32'h2308c; force soc.dbg_do = 32'h01079793; #1000;
force soc.dbg_adr = 32'h23090; force soc.dbg_do = 32'h0107d793; #1000;
force soc.dbg_adr = 32'h23094; force soc.dbg_do = 32'h0108d893; #1000;
force soc.dbg_adr = 32'h23098; force soc.dbg_do = 32'h418584b3; #1000;
force soc.dbg_adr = 32'h2309c; force soc.dbg_do = 32'h010bdb93; #1000;
force soc.dbg_adr = 32'h230a0; force soc.dbg_do = 32'h01095713; #1000;
force soc.dbg_adr = 32'h230a4; force soc.dbg_do = 32'h00078513; #1000;
force soc.dbg_adr = 32'h230a8; force soc.dbg_do = 32'h00088593; #1000;
force soc.dbg_adr = 32'h230ac; force soc.dbg_do = 32'h1a5000ef; #1000;
force soc.dbg_adr = 32'h230b0; force soc.dbg_do = 32'h00050813; #1000;
force soc.dbg_adr = 32'h230b4; force soc.dbg_do = 32'h00070593; #1000;
force soc.dbg_adr = 32'h230b8; force soc.dbg_do = 32'h00078513; #1000;
force soc.dbg_adr = 32'h230bc; force soc.dbg_do = 32'h00070793; #1000;
force soc.dbg_adr = 32'h230c0; force soc.dbg_do = 32'h191000ef; #1000;
force soc.dbg_adr = 32'h230c4; force soc.dbg_do = 32'h00050713; #1000;
force soc.dbg_adr = 32'h230c8; force soc.dbg_do = 32'h00088593; #1000;
force soc.dbg_adr = 32'h230cc; force soc.dbg_do = 32'h000b8513; #1000;
force soc.dbg_adr = 32'h230d0; force soc.dbg_do = 32'h181000ef; #1000;
force soc.dbg_adr = 32'h230d4; force soc.dbg_do = 32'h00050893; #1000;
force soc.dbg_adr = 32'h230d8; force soc.dbg_do = 32'h00078593; #1000;
force soc.dbg_adr = 32'h230dc; force soc.dbg_do = 32'h000b8513; #1000;
force soc.dbg_adr = 32'h230e0; force soc.dbg_do = 32'h171000ef; #1000;
force soc.dbg_adr = 32'h230e4; force soc.dbg_do = 32'h01085793; #1000;
force soc.dbg_adr = 32'h230e8; force soc.dbg_do = 32'h01170733; #1000;
force soc.dbg_adr = 32'h230ec; force soc.dbg_do = 32'h00e787b3; #1000;
force soc.dbg_adr = 32'h230f0; force soc.dbg_do = 32'h00050693; #1000;
force soc.dbg_adr = 32'h230f4; force soc.dbg_do = 32'h0117f663; #1000;
force soc.dbg_adr = 32'h230f8; force soc.dbg_do = 32'h00010737; #1000;
force soc.dbg_adr = 32'h230fc; force soc.dbg_do = 32'h00e506b3; #1000;
force soc.dbg_adr = 32'h23100; force soc.dbg_do = 32'h0107d713; #1000;
force soc.dbg_adr = 32'h23104; force soc.dbg_do = 32'h01081813; #1000;
force soc.dbg_adr = 32'h23108; force soc.dbg_do = 32'h01079793; #1000;
force soc.dbg_adr = 32'h2310c; force soc.dbg_do = 32'h01085813; #1000;
force soc.dbg_adr = 32'h23110; force soc.dbg_do = 32'h00d70733; #1000;
force soc.dbg_adr = 32'h23114; force soc.dbg_do = 32'h010787b3; #1000;
force soc.dbg_adr = 32'h23118; force soc.dbg_do = 32'h00e4e663; #1000;
force soc.dbg_adr = 32'h2311c; force soc.dbg_do = 32'h00e49e63; #1000;
force soc.dbg_adr = 32'h23120; force soc.dbg_do = 32'h00f9fc63; #1000;
force soc.dbg_adr = 32'h23124; force soc.dbg_do = 32'h41278933; #1000;
force soc.dbg_adr = 32'h23128; force soc.dbg_do = 32'h0127b6b3; #1000;
force soc.dbg_adr = 32'h2312c; force soc.dbg_do = 32'h016686b3; #1000;
force soc.dbg_adr = 32'h23130; force soc.dbg_do = 32'h00090793; #1000;
force soc.dbg_adr = 32'h23134; force soc.dbg_do = 32'h40d70733; #1000;
force soc.dbg_adr = 32'h23138; force soc.dbg_do = 32'h40f987b3; #1000;
force soc.dbg_adr = 32'h2313c; force soc.dbg_do = 32'h00f9b9b3; #1000;
force soc.dbg_adr = 32'h23140; force soc.dbg_do = 32'h40e485b3; #1000;
force soc.dbg_adr = 32'h23144; force soc.dbg_do = 32'h413585b3; #1000;
force soc.dbg_adr = 32'h23148; force soc.dbg_do = 32'h01559ab3; #1000;
force soc.dbg_adr = 32'h2314c; force soc.dbg_do = 32'h0147d7b3; #1000;
force soc.dbg_adr = 32'h23150; force soc.dbg_do = 32'h00fae533; #1000;
force soc.dbg_adr = 32'h23154; force soc.dbg_do = 32'h0145d5b3; #1000;
force soc.dbg_adr = 32'h23158; force soc.dbg_do = 32'hc71ff06f; #1000;
force soc.dbg_adr = 32'h2315c; force soc.dbg_do = 32'hfb010113; #1000;
force soc.dbg_adr = 32'h23160; force soc.dbg_do = 32'h03512a23; #1000;
force soc.dbg_adr = 32'h23164; force soc.dbg_do = 32'h0145da93; #1000;
force soc.dbg_adr = 32'h23168; force soc.dbg_do = 32'h04812423; #1000;
force soc.dbg_adr = 32'h2316c; force soc.dbg_do = 32'h03412c23; #1000;
force soc.dbg_adr = 32'h23170; force soc.dbg_do = 32'h03612823; #1000;
force soc.dbg_adr = 32'h23174; force soc.dbg_do = 32'h03812423; #1000;
force soc.dbg_adr = 32'h23178; force soc.dbg_do = 32'h03a12023; #1000;
force soc.dbg_adr = 32'h2317c; force soc.dbg_do = 32'h00c59413; #1000;
force soc.dbg_adr = 32'h23180; force soc.dbg_do = 32'h04112623; #1000;
force soc.dbg_adr = 32'h23184; force soc.dbg_do = 32'h04912223; #1000;
force soc.dbg_adr = 32'h23188; force soc.dbg_do = 32'h05212023; #1000;
force soc.dbg_adr = 32'h2318c; force soc.dbg_do = 32'h03312e23; #1000;
force soc.dbg_adr = 32'h23190; force soc.dbg_do = 32'h03712623; #1000;
force soc.dbg_adr = 32'h23194; force soc.dbg_do = 32'h03912223; #1000;
force soc.dbg_adr = 32'h23198; force soc.dbg_do = 32'h01b12e23; #1000;
force soc.dbg_adr = 32'h2319c; force soc.dbg_do = 32'h7ffafa93; #1000;
force soc.dbg_adr = 32'h231a0; force soc.dbg_do = 32'h00050a13; #1000;
force soc.dbg_adr = 32'h231a4; force soc.dbg_do = 32'h00060d13; #1000;
force soc.dbg_adr = 32'h231a8; force soc.dbg_do = 32'h00068c13; #1000;
force soc.dbg_adr = 32'h231ac; force soc.dbg_do = 32'h00c45413; #1000;
force soc.dbg_adr = 32'h231b0; force soc.dbg_do = 32'h01f5db13; #1000;
force soc.dbg_adr = 32'h231b4; force soc.dbg_do = 32'h0a0a8063; #1000;
force soc.dbg_adr = 32'h231b8; force soc.dbg_do = 32'h7ff00793; #1000;
force soc.dbg_adr = 32'h231bc; force soc.dbg_do = 32'h10fa8063; #1000;
force soc.dbg_adr = 32'h231c0; force soc.dbg_do = 32'h01d55b93; #1000;
force soc.dbg_adr = 32'h231c4; force soc.dbg_do = 32'h00341413; #1000;
force soc.dbg_adr = 32'h231c8; force soc.dbg_do = 32'h008bebb3; #1000;
force soc.dbg_adr = 32'h231cc; force soc.dbg_do = 32'h008007b7; #1000;
force soc.dbg_adr = 32'h231d0; force soc.dbg_do = 32'h00fbebb3; #1000;
force soc.dbg_adr = 32'h231d4; force soc.dbg_do = 32'h00351493; #1000;
force soc.dbg_adr = 32'h231d8; force soc.dbg_do = 32'hc01a8a93; #1000;
force soc.dbg_adr = 32'h231dc; force soc.dbg_do = 32'h00000c93; #1000;
force soc.dbg_adr = 32'h231e0; force soc.dbg_do = 32'h014c5713; #1000;
force soc.dbg_adr = 32'h231e4; force soc.dbg_do = 32'h00cc1413; #1000;
force soc.dbg_adr = 32'h231e8; force soc.dbg_do = 32'h7ff77713; #1000;
force soc.dbg_adr = 32'h231ec; force soc.dbg_do = 32'h00c45413; #1000;
force soc.dbg_adr = 32'h231f0; force soc.dbg_do = 32'h01fc5c13; #1000;
force soc.dbg_adr = 32'h231f4; force soc.dbg_do = 32'h0e070e63; #1000;
force soc.dbg_adr = 32'h231f8; force soc.dbg_do = 32'h7ff00793; #1000;
force soc.dbg_adr = 32'h231fc; force soc.dbg_do = 32'h16f70263; #1000;
force soc.dbg_adr = 32'h23200; force soc.dbg_do = 32'h00341413; #1000;
force soc.dbg_adr = 32'h23204; force soc.dbg_do = 32'h01dd5793; #1000;
force soc.dbg_adr = 32'h23208; force soc.dbg_do = 32'h0087e7b3; #1000;
force soc.dbg_adr = 32'h2320c; force soc.dbg_do = 32'h00800437; #1000;
force soc.dbg_adr = 32'h23210; force soc.dbg_do = 32'h0087e433; #1000;
force soc.dbg_adr = 32'h23214; force soc.dbg_do = 32'h003d1813; #1000;
force soc.dbg_adr = 32'h23218; force soc.dbg_do = 32'hc0170713; #1000;
force soc.dbg_adr = 32'h2321c; force soc.dbg_do = 32'h00000693; #1000;
force soc.dbg_adr = 32'h23220; force soc.dbg_do = 32'h002c9793; #1000;
force soc.dbg_adr = 32'h23224; force soc.dbg_do = 32'h00d7e7b3; #1000;
force soc.dbg_adr = 32'h23228; force soc.dbg_do = 32'h40ea8ab3; #1000;
force soc.dbg_adr = 32'h2322c; force soc.dbg_do = 32'hfff78793; #1000;
force soc.dbg_adr = 32'h23230; force soc.dbg_do = 32'h00e00713; #1000;
force soc.dbg_adr = 32'h23234; force soc.dbg_do = 32'h018b4a33; #1000;
force soc.dbg_adr = 32'h23238; force soc.dbg_do = 32'h14f76c63; #1000;
force soc.dbg_adr = 32'h2323c; force soc.dbg_do = 32'h00024737; #1000;
force soc.dbg_adr = 32'h23240; force soc.dbg_do = 32'h00279793; #1000;
force soc.dbg_adr = 32'h23244; force soc.dbg_do = 32'h1cc70713; #1000;
force soc.dbg_adr = 32'h23248; force soc.dbg_do = 32'h00e787b3; #1000;
force soc.dbg_adr = 32'h2324c; force soc.dbg_do = 32'h0007a783; #1000;
force soc.dbg_adr = 32'h23250; force soc.dbg_do = 32'h00078067; #1000;
force soc.dbg_adr = 32'h23254; force soc.dbg_do = 32'h00a46bb3; #1000;
force soc.dbg_adr = 32'h23258; force soc.dbg_do = 32'h060b8c63; #1000;
force soc.dbg_adr = 32'h2325c; force soc.dbg_do = 32'h02040e63; #1000;
force soc.dbg_adr = 32'h23260; force soc.dbg_do = 32'h00040513; #1000;
force soc.dbg_adr = 32'h23264; force soc.dbg_do = 32'h0c5000ef; #1000;
force soc.dbg_adr = 32'h23268; force soc.dbg_do = 32'hff550793; #1000;
force soc.dbg_adr = 32'h2326c; force soc.dbg_do = 32'h01d00b93; #1000;
force soc.dbg_adr = 32'h23270; force soc.dbg_do = 32'hff850713; #1000;
force soc.dbg_adr = 32'h23274; force soc.dbg_do = 32'h40fb8bb3; #1000;
force soc.dbg_adr = 32'h23278; force soc.dbg_do = 32'h00e41433; #1000;
force soc.dbg_adr = 32'h2327c; force soc.dbg_do = 32'h017a5bb3; #1000;
force soc.dbg_adr = 32'h23280; force soc.dbg_do = 32'h008bebb3; #1000;
force soc.dbg_adr = 32'h23284; force soc.dbg_do = 32'h00ea1433; #1000;
force soc.dbg_adr = 32'h23288; force soc.dbg_do = 32'hc0d00a93; #1000;
force soc.dbg_adr = 32'h2328c; force soc.dbg_do = 32'h40aa8ab3; #1000;
force soc.dbg_adr = 32'h23290; force soc.dbg_do = 32'h00040493; #1000;
force soc.dbg_adr = 32'h23294; force soc.dbg_do = 32'hf49ff06f; #1000;
force soc.dbg_adr = 32'h23298; force soc.dbg_do = 32'h091000ef; #1000;
force soc.dbg_adr = 32'h2329c; force soc.dbg_do = 32'h00050b93; #1000;
force soc.dbg_adr = 32'h232a0; force soc.dbg_do = 32'h015b8793; #1000;
force soc.dbg_adr = 32'h232a4; force soc.dbg_do = 32'h01c00713; #1000;
force soc.dbg_adr = 32'h232a8; force soc.dbg_do = 32'h02050513; #1000;
force soc.dbg_adr = 32'h232ac; force soc.dbg_do = 32'hfcf750e3; #1000;
force soc.dbg_adr = 32'h232b0; force soc.dbg_do = 32'hff8b8b93; #1000;
force soc.dbg_adr = 32'h232b4; force soc.dbg_do = 32'h017a1bb3; #1000;
force soc.dbg_adr = 32'h232b8; force soc.dbg_do = 32'hfd1ff06f; #1000;
force soc.dbg_adr = 32'h232bc; force soc.dbg_do = 32'h00a46bb3; #1000;
force soc.dbg_adr = 32'h232c0; force soc.dbg_do = 32'h020b9063; #1000;
force soc.dbg_adr = 32'h232c4; force soc.dbg_do = 32'h00000493; #1000;
force soc.dbg_adr = 32'h232c8; force soc.dbg_do = 32'h00200c93; #1000;
force soc.dbg_adr = 32'h232cc; force soc.dbg_do = 32'hf15ff06f; #1000;
force soc.dbg_adr = 32'h232d0; force soc.dbg_do = 32'h00000493; #1000;
force soc.dbg_adr = 32'h232d4; force soc.dbg_do = 32'h00000a93; #1000;
force soc.dbg_adr = 32'h232d8; force soc.dbg_do = 32'h00100c93; #1000;
force soc.dbg_adr = 32'h232dc; force soc.dbg_do = 32'hf05ff06f; #1000;
force soc.dbg_adr = 32'h232e0; force soc.dbg_do = 32'h00050493; #1000;
force soc.dbg_adr = 32'h232e4; force soc.dbg_do = 32'h00040b93; #1000;
force soc.dbg_adr = 32'h232e8; force soc.dbg_do = 32'h00300c93; #1000;
force soc.dbg_adr = 32'h232ec; force soc.dbg_do = 32'hef5ff06f; #1000;
force soc.dbg_adr = 32'h232f0; force soc.dbg_do = 32'h01a46833; #1000;
force soc.dbg_adr = 32'h232f4; force soc.dbg_do = 32'h08080063; #1000;
force soc.dbg_adr = 32'h232f8; force soc.dbg_do = 32'h04040063; #1000;
force soc.dbg_adr = 32'h232fc; force soc.dbg_do = 32'h00040513; #1000;
force soc.dbg_adr = 32'h23300; force soc.dbg_do = 32'h029000ef; #1000;
force soc.dbg_adr = 32'h23304; force soc.dbg_do = 32'hff550713; #1000;
force soc.dbg_adr = 32'h23308; force soc.dbg_do = 32'h01d00793; #1000;
force soc.dbg_adr = 32'h2330c; force soc.dbg_do = 32'hff850693; #1000;
force soc.dbg_adr = 32'h23310; force soc.dbg_do = 32'h40e787b3; #1000;
force soc.dbg_adr = 32'h23314; force soc.dbg_do = 32'h00d41433; #1000;
force soc.dbg_adr = 32'h23318; force soc.dbg_do = 32'h00fd57b3; #1000;
force soc.dbg_adr = 32'h2331c; force soc.dbg_do = 32'h0087e7b3; #1000;
force soc.dbg_adr = 32'h23320; force soc.dbg_do = 32'h00dd1433; #1000;
force soc.dbg_adr = 32'h23324; force soc.dbg_do = 32'hc0d00713; #1000;
force soc.dbg_adr = 32'h23328; force soc.dbg_do = 32'h00040813; #1000;
force soc.dbg_adr = 32'h2332c; force soc.dbg_do = 32'h40a70733; #1000;
force soc.dbg_adr = 32'h23330; force soc.dbg_do = 32'h00078413; #1000;
force soc.dbg_adr = 32'h23334; force soc.dbg_do = 32'hee9ff06f; #1000;
force soc.dbg_adr = 32'h23338; force soc.dbg_do = 32'h000d0513; #1000;
force soc.dbg_adr = 32'h2333c; force soc.dbg_do = 32'h7ec000ef; #1000;
force soc.dbg_adr = 32'h23340; force soc.dbg_do = 32'h00050793; #1000;
force soc.dbg_adr = 32'h23344; force soc.dbg_do = 32'h01578713; #1000;
force soc.dbg_adr = 32'h23348; force soc.dbg_do = 32'h01c00693; #1000;
force soc.dbg_adr = 32'h2334c; force soc.dbg_do = 32'h02050513; #1000;
force soc.dbg_adr = 32'h23350; force soc.dbg_do = 32'hfae6dce3; #1000;
force soc.dbg_adr = 32'h23354; force soc.dbg_do = 32'hff878793; #1000;
force soc.dbg_adr = 32'h23358; force soc.dbg_do = 32'h00fd17b3; #1000;
force soc.dbg_adr = 32'h2335c; force soc.dbg_do = 32'hfc9ff06f; #1000;
force soc.dbg_adr = 32'h23360; force soc.dbg_do = 32'h01a46833; #1000;
force soc.dbg_adr = 32'h23364; force soc.dbg_do = 32'h02081063; #1000;
force soc.dbg_adr = 32'h23368; force soc.dbg_do = 32'h00000413; #1000;
force soc.dbg_adr = 32'h2336c; force soc.dbg_do = 32'h00200693; #1000;
force soc.dbg_adr = 32'h23370; force soc.dbg_do = 32'heb1ff06f; #1000;
force soc.dbg_adr = 32'h23374; force soc.dbg_do = 32'h00000413; #1000;
force soc.dbg_adr = 32'h23378; force soc.dbg_do = 32'h00000713; #1000;
force soc.dbg_adr = 32'h2337c; force soc.dbg_do = 32'h00100693; #1000;
force soc.dbg_adr = 32'h23380; force soc.dbg_do = 32'hea1ff06f; #1000;
force soc.dbg_adr = 32'h23384; force soc.dbg_do = 32'h000d0813; #1000;
force soc.dbg_adr = 32'h23388; force soc.dbg_do = 32'h00300693; #1000;
force soc.dbg_adr = 32'h2338c; force soc.dbg_do = 32'he95ff06f; #1000;
force soc.dbg_adr = 32'h23390; force soc.dbg_do = 32'h01746663; #1000;
force soc.dbg_adr = 32'h23394; force soc.dbg_do = 32'h448b9e63; #1000;
force soc.dbg_adr = 32'h23398; force soc.dbg_do = 32'h4504ec63; #1000;
force soc.dbg_adr = 32'h2339c; force soc.dbg_do = 32'h01fb9713; #1000;
force soc.dbg_adr = 32'h233a0; force soc.dbg_do = 32'h0014d793; #1000;
force soc.dbg_adr = 32'h233a4; force soc.dbg_do = 32'h01f49c93; #1000;
force soc.dbg_adr = 32'h233a8; force soc.dbg_do = 32'h001bdb93; #1000;
force soc.dbg_adr = 32'h233ac; force soc.dbg_do = 32'h00f764b3; #1000;
force soc.dbg_adr = 32'h233b0; force soc.dbg_do = 32'h00841413; #1000;
force soc.dbg_adr = 32'h233b4; force soc.dbg_do = 32'h01045793; #1000;
force soc.dbg_adr = 32'h233b8; force soc.dbg_do = 32'h01885d93; #1000;
force soc.dbg_adr = 32'h233bc; force soc.dbg_do = 32'h00f12423; #1000;
force soc.dbg_adr = 32'h233c0; force soc.dbg_do = 32'h008dedb3; #1000;
force soc.dbg_adr = 32'h233c4; force soc.dbg_do = 32'h00812583; #1000;
force soc.dbg_adr = 32'h233c8; force soc.dbg_do = 32'h010d9793; #1000;
force soc.dbg_adr = 32'h233cc; force soc.dbg_do = 32'h0107d793; #1000;
force soc.dbg_adr = 32'h233d0; force soc.dbg_do = 32'h000b8513; #1000;
force soc.dbg_adr = 32'h233d4; force soc.dbg_do = 32'h00f12623; #1000;
force soc.dbg_adr = 32'h233d8; force soc.dbg_do = 32'h00881b13; #1000;
force soc.dbg_adr = 32'h233dc; force soc.dbg_do = 32'h6a0000ef; #1000;
force soc.dbg_adr = 32'h233e0; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h233e4; force soc.dbg_do = 32'h00050c13; #1000;
force soc.dbg_adr = 32'h233e8; force soc.dbg_do = 32'h010d9513; #1000;
force soc.dbg_adr = 32'h233ec; force soc.dbg_do = 32'h01055513; #1000;
force soc.dbg_adr = 32'h233f0; force soc.dbg_do = 32'h660000ef; #1000;
force soc.dbg_adr = 32'h233f4; force soc.dbg_do = 32'h00812583; #1000;
force soc.dbg_adr = 32'h233f8; force soc.dbg_do = 32'h00050413; #1000;
force soc.dbg_adr = 32'h233fc; force soc.dbg_do = 32'h000b8513; #1000;
force soc.dbg_adr = 32'h23400; force soc.dbg_do = 32'h6c4000ef; #1000;
force soc.dbg_adr = 32'h23404; force soc.dbg_do = 32'h01051513; #1000;
force soc.dbg_adr = 32'h23408; force soc.dbg_do = 32'h0104d793; #1000;
force soc.dbg_adr = 32'h2340c; force soc.dbg_do = 32'h00a7e7b3; #1000;
force soc.dbg_adr = 32'h23410; force soc.dbg_do = 32'h000c0b93; #1000;
force soc.dbg_adr = 32'h23414; force soc.dbg_do = 32'h0087fe63; #1000;
force soc.dbg_adr = 32'h23418; force soc.dbg_do = 32'h00fd87b3; #1000;
force soc.dbg_adr = 32'h2341c; force soc.dbg_do = 32'hfffc0b93; #1000;
force soc.dbg_adr = 32'h23420; force soc.dbg_do = 32'h01b7e863; #1000;
force soc.dbg_adr = 32'h23424; force soc.dbg_do = 32'h0087f663; #1000;
force soc.dbg_adr = 32'h23428; force soc.dbg_do = 32'hffec0b93; #1000;
force soc.dbg_adr = 32'h2342c; force soc.dbg_do = 32'h01b787b3; #1000;
force soc.dbg_adr = 32'h23430; force soc.dbg_do = 32'h00812583; #1000;
force soc.dbg_adr = 32'h23434; force soc.dbg_do = 32'h40878433; #1000;
force soc.dbg_adr = 32'h23438; force soc.dbg_do = 32'h00040513; #1000;
force soc.dbg_adr = 32'h2343c; force soc.dbg_do = 32'h640000ef; #1000;
force soc.dbg_adr = 32'h23440; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h23444; force soc.dbg_do = 32'h00050d13; #1000;
force soc.dbg_adr = 32'h23448; force soc.dbg_do = 32'h010d9513; #1000;
force soc.dbg_adr = 32'h2344c; force soc.dbg_do = 32'h01055513; #1000;
force soc.dbg_adr = 32'h23450; force soc.dbg_do = 32'h600000ef; #1000;
force soc.dbg_adr = 32'h23454; force soc.dbg_do = 32'h00812583; #1000;
force soc.dbg_adr = 32'h23458; force soc.dbg_do = 32'h00050c13; #1000;
force soc.dbg_adr = 32'h2345c; force soc.dbg_do = 32'h00040513; #1000;
force soc.dbg_adr = 32'h23460; force soc.dbg_do = 32'h664000ef; #1000;
force soc.dbg_adr = 32'h23464; force soc.dbg_do = 32'h01049493; #1000;
force soc.dbg_adr = 32'h23468; force soc.dbg_do = 32'h01051513; #1000;
force soc.dbg_adr = 32'h2346c; force soc.dbg_do = 32'h0104d493; #1000;
force soc.dbg_adr = 32'h23470; force soc.dbg_do = 32'h00a4e4b3; #1000;
force soc.dbg_adr = 32'h23474; force soc.dbg_do = 32'h000d0793; #1000;
force soc.dbg_adr = 32'h23478; force soc.dbg_do = 32'h0184fe63; #1000;
force soc.dbg_adr = 32'h2347c; force soc.dbg_do = 32'h009d84b3; #1000;
force soc.dbg_adr = 32'h23480; force soc.dbg_do = 32'hfffd0793; #1000;
force soc.dbg_adr = 32'h23484; force soc.dbg_do = 32'h01b4e863; #1000;
force soc.dbg_adr = 32'h23488; force soc.dbg_do = 32'h0184f663; #1000;
force soc.dbg_adr = 32'h2348c; force soc.dbg_do = 32'hffed0793; #1000;
force soc.dbg_adr = 32'h23490; force soc.dbg_do = 32'h01b484b3; #1000;
force soc.dbg_adr = 32'h23494; force soc.dbg_do = 32'h010b9813; #1000;
force soc.dbg_adr = 32'h23498; force soc.dbg_do = 32'h00f86833; #1000;
force soc.dbg_adr = 32'h2349c; force soc.dbg_do = 32'h01081793; #1000;
force soc.dbg_adr = 32'h234a0; force soc.dbg_do = 32'h010b1713; #1000;
force soc.dbg_adr = 32'h234a4; force soc.dbg_do = 32'h01075713; #1000;
force soc.dbg_adr = 32'h234a8; force soc.dbg_do = 32'h0107d793; #1000;
force soc.dbg_adr = 32'h234ac; force soc.dbg_do = 32'h418484b3; #1000;
force soc.dbg_adr = 32'h234b0; force soc.dbg_do = 32'h01085e93; #1000;
force soc.dbg_adr = 32'h234b4; force soc.dbg_do = 32'h00078513; #1000;
force soc.dbg_adr = 32'h234b8; force soc.dbg_do = 32'h00e12623; #1000;
force soc.dbg_adr = 32'h234bc; force soc.dbg_do = 32'h00070593; #1000;
force soc.dbg_adr = 32'h234c0; force soc.dbg_do = 32'h590000ef; #1000;
force soc.dbg_adr = 32'h234c4; force soc.dbg_do = 32'h00050313; #1000;
force soc.dbg_adr = 32'h234c8; force soc.dbg_do = 32'h010b5593; #1000;
force soc.dbg_adr = 32'h234cc; force soc.dbg_do = 32'h00078513; #1000;
force soc.dbg_adr = 32'h234d0; force soc.dbg_do = 32'h580000ef; #1000;
force soc.dbg_adr = 32'h234d4; force soc.dbg_do = 32'h00050793; #1000;
force soc.dbg_adr = 32'h234d8; force soc.dbg_do = 32'h00070593; #1000;
force soc.dbg_adr = 32'h234dc; force soc.dbg_do = 32'h000e8513; #1000;
force soc.dbg_adr = 32'h234e0; force soc.dbg_do = 32'h570000ef; #1000;
force soc.dbg_adr = 32'h234e4; force soc.dbg_do = 32'h00050e13; #1000;
force soc.dbg_adr = 32'h234e8; force soc.dbg_do = 32'h010b5593; #1000;
force soc.dbg_adr = 32'h234ec; force soc.dbg_do = 32'h000e8513; #1000;
force soc.dbg_adr = 32'h234f0; force soc.dbg_do = 32'h560000ef; #1000;
force soc.dbg_adr = 32'h234f4; force soc.dbg_do = 32'h01035d13; #1000;
force soc.dbg_adr = 32'h234f8; force soc.dbg_do = 32'h01c787b3; #1000;
force soc.dbg_adr = 32'h234fc; force soc.dbg_do = 32'h00fd0d33; #1000;
force soc.dbg_adr = 32'h23500; force soc.dbg_do = 32'h00050693; #1000;
force soc.dbg_adr = 32'h23504; force soc.dbg_do = 32'h01cd7663; #1000;
force soc.dbg_adr = 32'h23508; force soc.dbg_do = 32'h000107b7; #1000;
force soc.dbg_adr = 32'h2350c; force soc.dbg_do = 32'h00f506b3; #1000;
force soc.dbg_adr = 32'h23510; force soc.dbg_do = 32'h010d5793; #1000;
force soc.dbg_adr = 32'h23514; force soc.dbg_do = 32'h01031313; #1000;
force soc.dbg_adr = 32'h23518; force soc.dbg_do = 32'h010d1d13; #1000;
force soc.dbg_adr = 32'h2351c; force soc.dbg_do = 32'h01035313; #1000;
force soc.dbg_adr = 32'h23520; force soc.dbg_do = 32'h00d787b3; #1000;
force soc.dbg_adr = 32'h23524; force soc.dbg_do = 32'h006d0d33; #1000;
force soc.dbg_adr = 32'h23528; force soc.dbg_do = 32'h00f4e863; #1000;
force soc.dbg_adr = 32'h2352c; force soc.dbg_do = 32'h00080413; #1000;
force soc.dbg_adr = 32'h23530; force soc.dbg_do = 32'h04f49863; #1000;
force soc.dbg_adr = 32'h23534; force soc.dbg_do = 32'h05acf663; #1000;
force soc.dbg_adr = 32'h23538; force soc.dbg_do = 32'h016c86b3; #1000;
force soc.dbg_adr = 32'h2353c; force soc.dbg_do = 32'h0196b633; #1000;
force soc.dbg_adr = 32'h23540; force soc.dbg_do = 32'h01b605b3; #1000;
force soc.dbg_adr = 32'h23544; force soc.dbg_do = 32'h00b484b3; #1000;
force soc.dbg_adr = 32'h23548; force soc.dbg_do = 32'hfff80413; #1000;
force soc.dbg_adr = 32'h2354c; force soc.dbg_do = 32'h00068c93; #1000;
force soc.dbg_adr = 32'h23550; force soc.dbg_do = 32'h009de663; #1000;
force soc.dbg_adr = 32'h23554; force soc.dbg_do = 32'h029d9663; #1000;
force soc.dbg_adr = 32'h23558; force soc.dbg_do = 32'h02061463; #1000;
force soc.dbg_adr = 32'h2355c; force soc.dbg_do = 32'h00f4e663; #1000;
force soc.dbg_adr = 32'h23560; force soc.dbg_do = 32'h02979063; #1000;
force soc.dbg_adr = 32'h23564; force soc.dbg_do = 32'h01a6fe63; #1000;
force soc.dbg_adr = 32'h23568; force soc.dbg_do = 32'h00db06b3; #1000;
force soc.dbg_adr = 32'h2356c; force soc.dbg_do = 32'h00068c93; #1000;
force soc.dbg_adr = 32'h23570; force soc.dbg_do = 32'h0166b6b3; #1000;
force soc.dbg_adr = 32'h23574; force soc.dbg_do = 32'h01b686b3; #1000;
force soc.dbg_adr = 32'h23578; force soc.dbg_do = 32'hffe80413; #1000;
force soc.dbg_adr = 32'h2357c; force soc.dbg_do = 32'h00d484b3; #1000;
force soc.dbg_adr = 32'h23580; force soc.dbg_do = 32'h41ac8d33; #1000;
force soc.dbg_adr = 32'h23584; force soc.dbg_do = 32'h40f484b3; #1000;
force soc.dbg_adr = 32'h23588; force soc.dbg_do = 32'h01acb8b3; #1000;
force soc.dbg_adr = 32'h2358c; force soc.dbg_do = 32'h411484b3; #1000;
force soc.dbg_adr = 32'h23590; force soc.dbg_do = 32'hfff00813; #1000;
force soc.dbg_adr = 32'h23594; force soc.dbg_do = 32'h1a9d8263; #1000;
force soc.dbg_adr = 32'h23598; force soc.dbg_do = 32'h00812583; #1000;
force soc.dbg_adr = 32'h2359c; force soc.dbg_do = 32'h00048513; #1000;
force soc.dbg_adr = 32'h235a0; force soc.dbg_do = 32'h4dc000ef; #1000;
force soc.dbg_adr = 32'h235a4; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h235a8; force soc.dbg_do = 32'h00050c13; #1000;
force soc.dbg_adr = 32'h235ac; force soc.dbg_do = 32'h010d9513; #1000;
force soc.dbg_adr = 32'h235b0; force soc.dbg_do = 32'h01055513; #1000;
force soc.dbg_adr = 32'h235b4; force soc.dbg_do = 32'h49c000ef; #1000;
force soc.dbg_adr = 32'h235b8; force soc.dbg_do = 32'h00812583; #1000;
force soc.dbg_adr = 32'h235bc; force soc.dbg_do = 32'h00050b93; #1000;
force soc.dbg_adr = 32'h235c0; force soc.dbg_do = 32'h00048513; #1000;
force soc.dbg_adr = 32'h235c4; force soc.dbg_do = 32'h500000ef; #1000;
force soc.dbg_adr = 32'h235c8; force soc.dbg_do = 32'h01051513; #1000;
force soc.dbg_adr = 32'h235cc; force soc.dbg_do = 32'h010d5793; #1000;
force soc.dbg_adr = 32'h235d0; force soc.dbg_do = 32'h00a7e7b3; #1000;
force soc.dbg_adr = 32'h235d4; force soc.dbg_do = 32'h000c0493; #1000;
force soc.dbg_adr = 32'h235d8; force soc.dbg_do = 32'h0177fe63; #1000;
force soc.dbg_adr = 32'h235dc; force soc.dbg_do = 32'h00fd87b3; #1000;
force soc.dbg_adr = 32'h235e0; force soc.dbg_do = 32'hfffc0493; #1000;
force soc.dbg_adr = 32'h235e4; force soc.dbg_do = 32'h01b7e863; #1000;
force soc.dbg_adr = 32'h235e8; force soc.dbg_do = 32'h0177f663; #1000;
force soc.dbg_adr = 32'h235ec; force soc.dbg_do = 32'hffec0493; #1000;
force soc.dbg_adr = 32'h235f0; force soc.dbg_do = 32'h01b787b3; #1000;
force soc.dbg_adr = 32'h235f4; force soc.dbg_do = 32'h00812583; #1000;
force soc.dbg_adr = 32'h235f8; force soc.dbg_do = 32'h41778c33; #1000;
force soc.dbg_adr = 32'h235fc; force soc.dbg_do = 32'h000c0513; #1000;
force soc.dbg_adr = 32'h23600; force soc.dbg_do = 32'h47c000ef; #1000;
force soc.dbg_adr = 32'h23604; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h23608; force soc.dbg_do = 32'h00050b93; #1000;
force soc.dbg_adr = 32'h2360c; force soc.dbg_do = 32'h010d9513; #1000;
force soc.dbg_adr = 32'h23610; force soc.dbg_do = 32'h01055513; #1000;
force soc.dbg_adr = 32'h23614; force soc.dbg_do = 32'h43c000ef; #1000;
force soc.dbg_adr = 32'h23618; force soc.dbg_do = 32'h00812583; #1000;
force soc.dbg_adr = 32'h2361c; force soc.dbg_do = 32'h00050c93; #1000;
force soc.dbg_adr = 32'h23620; force soc.dbg_do = 32'h000c0513; #1000;
force soc.dbg_adr = 32'h23624; force soc.dbg_do = 32'h4a0000ef; #1000;
force soc.dbg_adr = 32'h23628; force soc.dbg_do = 32'h010d1793; #1000;
force soc.dbg_adr = 32'h2362c; force soc.dbg_do = 32'h01051513; #1000;
force soc.dbg_adr = 32'h23630; force soc.dbg_do = 32'h0107d793; #1000;
force soc.dbg_adr = 32'h23634; force soc.dbg_do = 32'h00a7e7b3; #1000;
force soc.dbg_adr = 32'h23638; force soc.dbg_do = 32'h000b8613; #1000;
force soc.dbg_adr = 32'h2363c; force soc.dbg_do = 32'h0197fe63; #1000;
force soc.dbg_adr = 32'h23640; force soc.dbg_do = 32'h00fd87b3; #1000;
force soc.dbg_adr = 32'h23644; force soc.dbg_do = 32'hfffb8613; #1000;
force soc.dbg_adr = 32'h23648; force soc.dbg_do = 32'h01b7e863; #1000;
force soc.dbg_adr = 32'h2364c; force soc.dbg_do = 32'h0197f663; #1000;
force soc.dbg_adr = 32'h23650; force soc.dbg_do = 32'hffeb8613; #1000;
force soc.dbg_adr = 32'h23654; force soc.dbg_do = 32'h01b787b3; #1000;
force soc.dbg_adr = 32'h23658; force soc.dbg_do = 32'h01049893; #1000;
force soc.dbg_adr = 32'h2365c; force soc.dbg_do = 32'h00c8e8b3; #1000;
force soc.dbg_adr = 32'h23660; force soc.dbg_do = 32'h01089313; #1000;
force soc.dbg_adr = 32'h23664; force soc.dbg_do = 32'h01035313; #1000;
force soc.dbg_adr = 32'h23668; force soc.dbg_do = 32'h010b1593; #1000;
force soc.dbg_adr = 32'h2366c; force soc.dbg_do = 32'h419787b3; #1000;
force soc.dbg_adr = 32'h23670; force soc.dbg_do = 32'h0108de93; #1000;
force soc.dbg_adr = 32'h23674; force soc.dbg_do = 32'h00030513; #1000;
force soc.dbg_adr = 32'h23678; force soc.dbg_do = 32'h0105d593; #1000;
force soc.dbg_adr = 32'h2367c; force soc.dbg_do = 32'h3d4000ef; #1000;
force soc.dbg_adr = 32'h23680; force soc.dbg_do = 32'h00050813; #1000;
force soc.dbg_adr = 32'h23684; force soc.dbg_do = 32'h010b5593; #1000;
force soc.dbg_adr = 32'h23688; force soc.dbg_do = 32'h00030513; #1000;
force soc.dbg_adr = 32'h2368c; force soc.dbg_do = 32'h3c4000ef; #1000;
force soc.dbg_adr = 32'h23690; force soc.dbg_do = 32'h010b1593; #1000;
force soc.dbg_adr = 32'h23694; force soc.dbg_do = 32'h00050313; #1000;
force soc.dbg_adr = 32'h23698; force soc.dbg_do = 32'h0105d593; #1000;
force soc.dbg_adr = 32'h2369c; force soc.dbg_do = 32'h000e8513; #1000;
force soc.dbg_adr = 32'h236a0; force soc.dbg_do = 32'h3b0000ef; #1000;
force soc.dbg_adr = 32'h236a4; force soc.dbg_do = 32'h00050e13; #1000;
force soc.dbg_adr = 32'h236a8; force soc.dbg_do = 32'h010b5593; #1000;
force soc.dbg_adr = 32'h236ac; force soc.dbg_do = 32'h000e8513; #1000;
force soc.dbg_adr = 32'h236b0; force soc.dbg_do = 32'h3a0000ef; #1000;
force soc.dbg_adr = 32'h236b4; force soc.dbg_do = 32'h01085693; #1000;
force soc.dbg_adr = 32'h236b8; force soc.dbg_do = 32'h01c30333; #1000;
force soc.dbg_adr = 32'h236bc; force soc.dbg_do = 32'h006686b3; #1000;
force soc.dbg_adr = 32'h236c0; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h236c4; force soc.dbg_do = 32'h01c6f663; #1000;
force soc.dbg_adr = 32'h236c8; force soc.dbg_do = 32'h00010637; #1000;
force soc.dbg_adr = 32'h236cc; force soc.dbg_do = 32'h00c505b3; #1000;
force soc.dbg_adr = 32'h236d0; force soc.dbg_do = 32'h0106d613; #1000;
force soc.dbg_adr = 32'h236d4; force soc.dbg_do = 32'h01081813; #1000;
force soc.dbg_adr = 32'h236d8; force soc.dbg_do = 32'h01069693; #1000;
force soc.dbg_adr = 32'h236dc; force soc.dbg_do = 32'h01085813; #1000;
force soc.dbg_adr = 32'h236e0; force soc.dbg_do = 32'h00b60633; #1000;
force soc.dbg_adr = 32'h236e4; force soc.dbg_do = 32'h010686b3; #1000;
force soc.dbg_adr = 32'h236e8; force soc.dbg_do = 32'h00c7e863; #1000;
force soc.dbg_adr = 32'h236ec; force soc.dbg_do = 32'h00088813; #1000;
force soc.dbg_adr = 32'h236f0; force soc.dbg_do = 32'h04c79263; #1000;
force soc.dbg_adr = 32'h236f4; force soc.dbg_do = 32'h04068263; #1000;
force soc.dbg_adr = 32'h236f8; force soc.dbg_do = 32'h00fd87b3; #1000;
force soc.dbg_adr = 32'h236fc; force soc.dbg_do = 32'hfff88813; #1000;
force soc.dbg_adr = 32'h23700; force soc.dbg_do = 32'h00078593; #1000;
force soc.dbg_adr = 32'h23704; force soc.dbg_do = 32'h03b7e463; #1000;
force soc.dbg_adr = 32'h23708; force soc.dbg_do = 32'h00c7e663; #1000;
force soc.dbg_adr = 32'h2370c; force soc.dbg_do = 32'h02c79463; #1000;
force soc.dbg_adr = 32'h23710; force soc.dbg_do = 32'h02db7063; #1000;
force soc.dbg_adr = 32'h23714; force soc.dbg_do = 32'h001b1513; #1000;
force soc.dbg_adr = 32'h23718; force soc.dbg_do = 32'h016535b3; #1000;
force soc.dbg_adr = 32'h2371c; force soc.dbg_do = 32'h01b585b3; #1000;
force soc.dbg_adr = 32'h23720; force soc.dbg_do = 32'hffe88813; #1000;
force soc.dbg_adr = 32'h23724; force soc.dbg_do = 32'h00b785b3; #1000;
force soc.dbg_adr = 32'h23728; force soc.dbg_do = 32'h00050b13; #1000;
force soc.dbg_adr = 32'h2372c; force soc.dbg_do = 32'h00c59463; #1000;
force soc.dbg_adr = 32'h23730; force soc.dbg_do = 32'h01668463; #1000;
force soc.dbg_adr = 32'h23734; force soc.dbg_do = 32'h00186813; #1000;
force soc.dbg_adr = 32'h23738; force soc.dbg_do = 32'h3ffa8793; #1000;
force soc.dbg_adr = 32'h2373c; force soc.dbg_do = 32'h0ef05e63; #1000;
force soc.dbg_adr = 32'h23740; force soc.dbg_do = 32'h00787713; #1000;
force soc.dbg_adr = 32'h23744; force soc.dbg_do = 32'h02070063; #1000;
force soc.dbg_adr = 32'h23748; force soc.dbg_do = 32'h00f87713; #1000;
force soc.dbg_adr = 32'h2374c; force soc.dbg_do = 32'h00400693; #1000;
force soc.dbg_adr = 32'h23750; force soc.dbg_do = 32'h00d70a63; #1000;
force soc.dbg_adr = 32'h23754; force soc.dbg_do = 32'h00d80733; #1000;
force soc.dbg_adr = 32'h23758; force soc.dbg_do = 32'h010736b3; #1000;
force soc.dbg_adr = 32'h2375c; force soc.dbg_do = 32'h00d40433; #1000;
force soc.dbg_adr = 32'h23760; force soc.dbg_do = 32'h00070813; #1000;
force soc.dbg_adr = 32'h23764; force soc.dbg_do = 32'h00741713; #1000;
force soc.dbg_adr = 32'h23768; force soc.dbg_do = 32'h00075a63; #1000;
force soc.dbg_adr = 32'h2376c; force soc.dbg_do = 32'hff0007b7; #1000;
force soc.dbg_adr = 32'h23770; force soc.dbg_do = 32'hfff78793; #1000;
force soc.dbg_adr = 32'h23774; force soc.dbg_do = 32'h00f47433; #1000;
force soc.dbg_adr = 32'h23778; force soc.dbg_do = 32'h400a8793; #1000;
force soc.dbg_adr = 32'h2377c; force soc.dbg_do = 32'h7fe00713; #1000;
force soc.dbg_adr = 32'h23780; force soc.dbg_do = 32'h18f74063; #1000;
force soc.dbg_adr = 32'h23784; force soc.dbg_do = 32'h01d41713; #1000;
force soc.dbg_adr = 32'h23788; force soc.dbg_do = 32'h00385813; #1000;
force soc.dbg_adr = 32'h2378c; force soc.dbg_do = 32'h01076833; #1000;
force soc.dbg_adr = 32'h23790; force soc.dbg_do = 32'h00345413; #1000;
force soc.dbg_adr = 32'h23794; force soc.dbg_do = 32'h00c41413; #1000;
force soc.dbg_adr = 32'h23798; force soc.dbg_do = 32'h00c45413; #1000;
force soc.dbg_adr = 32'h2379c; force soc.dbg_do = 32'h01479793; #1000;
force soc.dbg_adr = 32'h237a0; force soc.dbg_do = 32'h04c12083; #1000;
force soc.dbg_adr = 32'h237a4; force soc.dbg_do = 32'h0087e7b3; #1000;
force soc.dbg_adr = 32'h237a8; force soc.dbg_do = 32'h04812403; #1000;
force soc.dbg_adr = 32'h237ac; force soc.dbg_do = 32'h01fa1a13; #1000;
force soc.dbg_adr = 32'h237b0; force soc.dbg_do = 32'h0147e733; #1000;
force soc.dbg_adr = 32'h237b4; force soc.dbg_do = 32'h04412483; #1000;
force soc.dbg_adr = 32'h237b8; force soc.dbg_do = 32'h04012903; #1000;
force soc.dbg_adr = 32'h237bc; force soc.dbg_do = 32'h03c12983; #1000;
force soc.dbg_adr = 32'h237c0; force soc.dbg_do = 32'h03812a03; #1000;
force soc.dbg_adr = 32'h237c4; force soc.dbg_do = 32'h03412a83; #1000;
force soc.dbg_adr = 32'h237c8; force soc.dbg_do = 32'h03012b03; #1000;
force soc.dbg_adr = 32'h237cc; force soc.dbg_do = 32'h02c12b83; #1000;
force soc.dbg_adr = 32'h237d0; force soc.dbg_do = 32'h02812c03; #1000;
force soc.dbg_adr = 32'h237d4; force soc.dbg_do = 32'h02412c83; #1000;
force soc.dbg_adr = 32'h237d8; force soc.dbg_do = 32'h02012d03; #1000;
force soc.dbg_adr = 32'h237dc; force soc.dbg_do = 32'h01c12d83; #1000;
force soc.dbg_adr = 32'h237e0; force soc.dbg_do = 32'h00080513; #1000;
force soc.dbg_adr = 32'h237e4; force soc.dbg_do = 32'h00070593; #1000;
force soc.dbg_adr = 32'h237e8; force soc.dbg_do = 32'h05010113; #1000;
force soc.dbg_adr = 32'h237ec; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h237f0; force soc.dbg_do = 32'hfffa8a93; #1000;
force soc.dbg_adr = 32'h237f4; force soc.dbg_do = 32'h00000c93; #1000;
force soc.dbg_adr = 32'h237f8; force soc.dbg_do = 32'hbb9ff06f; #1000;
force soc.dbg_adr = 32'h237fc; force soc.dbg_do = 32'h000c0a13; #1000;
force soc.dbg_adr = 32'h23800; force soc.dbg_do = 32'h00068c93; #1000;
force soc.dbg_adr = 32'h23804; force soc.dbg_do = 32'h00200793; #1000;
force soc.dbg_adr = 32'h23808; force soc.dbg_do = 32'h0efc8c63; #1000;
force soc.dbg_adr = 32'h2380c; force soc.dbg_do = 32'h00300793; #1000;
force soc.dbg_adr = 32'h23810; force soc.dbg_do = 32'h0cfc8e63; #1000;
force soc.dbg_adr = 32'h23814; force soc.dbg_do = 32'h00100793; #1000;
force soc.dbg_adr = 32'h23818; force soc.dbg_do = 32'hf2fc90e3; #1000;
force soc.dbg_adr = 32'h2381c; force soc.dbg_do = 32'h00000413; #1000;
force soc.dbg_adr = 32'h23820; force soc.dbg_do = 32'h00000813; #1000;
force soc.dbg_adr = 32'h23824; force soc.dbg_do = 32'h08c0006f; #1000;
force soc.dbg_adr = 32'h23828; force soc.dbg_do = 32'h000b0a13; #1000;
force soc.dbg_adr = 32'h2382c; force soc.dbg_do = 32'h000b8413; #1000;
force soc.dbg_adr = 32'h23830; force soc.dbg_do = 32'h00048813; #1000;
force soc.dbg_adr = 32'h23834; force soc.dbg_do = 32'hfd1ff06f; #1000;
force soc.dbg_adr = 32'h23838; force soc.dbg_do = 32'h00100693; #1000;
force soc.dbg_adr = 32'h2383c; force soc.dbg_do = 32'h00078c63; #1000;
force soc.dbg_adr = 32'h23840; force soc.dbg_do = 32'h40f686b3; #1000;
force soc.dbg_adr = 32'h23844; force soc.dbg_do = 32'h03800713; #1000;
force soc.dbg_adr = 32'h23848; force soc.dbg_do = 32'hfcd74ae3; #1000;
force soc.dbg_adr = 32'h2384c; force soc.dbg_do = 32'h01f00713; #1000;
force soc.dbg_adr = 32'h23850; force soc.dbg_do = 32'h06d74463; #1000;
force soc.dbg_adr = 32'h23854; force soc.dbg_do = 32'h41ea8a93; #1000;
force soc.dbg_adr = 32'h23858; force soc.dbg_do = 32'h00d857b3; #1000;
force soc.dbg_adr = 32'h2385c; force soc.dbg_do = 32'h01581833; #1000;
force soc.dbg_adr = 32'h23860; force soc.dbg_do = 32'h01003833; #1000;
force soc.dbg_adr = 32'h23864; force soc.dbg_do = 32'h01541ab3; #1000;
force soc.dbg_adr = 32'h23868; force soc.dbg_do = 32'h01586833; #1000;
force soc.dbg_adr = 32'h2386c; force soc.dbg_do = 32'h0107e7b3; #1000;
force soc.dbg_adr = 32'h23870; force soc.dbg_do = 32'h00d45433; #1000;
force soc.dbg_adr = 32'h23874; force soc.dbg_do = 32'h0077f713; #1000;
force soc.dbg_adr = 32'h23878; force soc.dbg_do = 32'h02070063; #1000;
force soc.dbg_adr = 32'h2387c; force soc.dbg_do = 32'h00f7f713; #1000;
force soc.dbg_adr = 32'h23880; force soc.dbg_do = 32'h00400693; #1000;
force soc.dbg_adr = 32'h23884; force soc.dbg_do = 32'h00d70a63; #1000;
force soc.dbg_adr = 32'h23888; force soc.dbg_do = 32'h00d78733; #1000;
force soc.dbg_adr = 32'h2388c; force soc.dbg_do = 32'h00f736b3; #1000;
force soc.dbg_adr = 32'h23890; force soc.dbg_do = 32'h00d40433; #1000;
force soc.dbg_adr = 32'h23894; force soc.dbg_do = 32'h00070793; #1000;
force soc.dbg_adr = 32'h23898; force soc.dbg_do = 32'h00841713; #1000;
force soc.dbg_adr = 32'h2389c; force soc.dbg_do = 32'h06074a63; #1000;
force soc.dbg_adr = 32'h238a0; force soc.dbg_do = 32'h01d41813; #1000;
force soc.dbg_adr = 32'h238a4; force soc.dbg_do = 32'h0037d793; #1000;
force soc.dbg_adr = 32'h238a8; force soc.dbg_do = 32'h00f86833; #1000;
force soc.dbg_adr = 32'h238ac; force soc.dbg_do = 32'h00345413; #1000;
force soc.dbg_adr = 32'h238b0; force soc.dbg_do = 32'h00000793; #1000;
force soc.dbg_adr = 32'h238b4; force soc.dbg_do = 32'hee1ff06f; #1000;
force soc.dbg_adr = 32'h238b8; force soc.dbg_do = 32'hfe100713; #1000;
force soc.dbg_adr = 32'h238bc; force soc.dbg_do = 32'h40f707b3; #1000;
force soc.dbg_adr = 32'h238c0; force soc.dbg_do = 32'h02000613; #1000;
force soc.dbg_adr = 32'h238c4; force soc.dbg_do = 32'h00f457b3; #1000;
force soc.dbg_adr = 32'h238c8; force soc.dbg_do = 32'h00000713; #1000;
force soc.dbg_adr = 32'h238cc; force soc.dbg_do = 32'h00c68663; #1000;
force soc.dbg_adr = 32'h238d0; force soc.dbg_do = 32'h43ea8a93; #1000;
force soc.dbg_adr = 32'h238d4; force soc.dbg_do = 32'h01541733; #1000;
force soc.dbg_adr = 32'h238d8; force soc.dbg_do = 32'h01076733; #1000;
force soc.dbg_adr = 32'h238dc; force soc.dbg_do = 32'h00e03733; #1000;
force soc.dbg_adr = 32'h238e0; force soc.dbg_do = 32'h00e7e7b3; #1000;
force soc.dbg_adr = 32'h238e4; force soc.dbg_do = 32'h00000413; #1000;
force soc.dbg_adr = 32'h238e8; force soc.dbg_do = 32'hf8dff06f; #1000;
force soc.dbg_adr = 32'h238ec; force soc.dbg_do = 32'h00080437; #1000;
force soc.dbg_adr = 32'h238f0; force soc.dbg_do = 32'h00000813; #1000;
force soc.dbg_adr = 32'h238f4; force soc.dbg_do = 32'h7ff00793; #1000;
force soc.dbg_adr = 32'h238f8; force soc.dbg_do = 32'h00000a13; #1000;
force soc.dbg_adr = 32'h238fc; force soc.dbg_do = 32'he99ff06f; #1000;
force soc.dbg_adr = 32'h23900; force soc.dbg_do = 32'h00000413; #1000;
force soc.dbg_adr = 32'h23904; force soc.dbg_do = 32'h00000813; #1000;
force soc.dbg_adr = 32'h23908; force soc.dbg_do = 32'h7ff00793; #1000;
force soc.dbg_adr = 32'h2390c; force soc.dbg_do = 32'he89ff06f; #1000;
force soc.dbg_adr = 32'h23910; force soc.dbg_do = 32'h00000413; #1000;
force soc.dbg_adr = 32'h23914; force soc.dbg_do = 32'h00000813; #1000;
force soc.dbg_adr = 32'h23918; force soc.dbg_do = 32'h00100793; #1000;
force soc.dbg_adr = 32'h2391c; force soc.dbg_do = 32'he79ff06f; #1000;
force soc.dbg_adr = 32'h23920; force soc.dbg_do = 32'h0145d713; #1000;
force soc.dbg_adr = 32'h23924; force soc.dbg_do = 32'h00100837; #1000;
force soc.dbg_adr = 32'h23928; force soc.dbg_do = 32'hfff80793; #1000;
force soc.dbg_adr = 32'h2392c; force soc.dbg_do = 32'h7ff77713; #1000;
force soc.dbg_adr = 32'h23930; force soc.dbg_do = 32'h3fe00613; #1000;
force soc.dbg_adr = 32'h23934; force soc.dbg_do = 32'h00b7f7b3; #1000;
force soc.dbg_adr = 32'h23938; force soc.dbg_do = 32'h00050693; #1000;
force soc.dbg_adr = 32'h2393c; force soc.dbg_do = 32'h01f5d593; #1000;
force soc.dbg_adr = 32'h23940; force soc.dbg_do = 32'h04e65a63; #1000;
force soc.dbg_adr = 32'h23944; force soc.dbg_do = 32'h41f00613; #1000;
force soc.dbg_adr = 32'h23948; force soc.dbg_do = 32'h40b60633; #1000;
force soc.dbg_adr = 32'h2394c; force soc.dbg_do = 32'hfff58513; #1000;
force soc.dbg_adr = 32'h23950; force soc.dbg_do = 32'h04c75463; #1000;
force soc.dbg_adr = 32'h23954; force soc.dbg_do = 32'h00000513; #1000;
force soc.dbg_adr = 32'h23958; force soc.dbg_do = 32'h04059063; #1000;
force soc.dbg_adr = 32'h2395c; force soc.dbg_do = 32'h43300613; #1000;
force soc.dbg_adr = 32'h23960; force soc.dbg_do = 32'h40e60633; #1000;
force soc.dbg_adr = 32'h23964; force soc.dbg_do = 32'h01f00593; #1000;
force soc.dbg_adr = 32'h23968; force soc.dbg_do = 32'h0107e7b3; #1000;
force soc.dbg_adr = 32'h2396c; force soc.dbg_do = 32'h00c5cc63; #1000;
force soc.dbg_adr = 32'h23970; force soc.dbg_do = 32'hbed70713; #1000;
force soc.dbg_adr = 32'h23974; force soc.dbg_do = 32'h00e797b3; #1000;
force soc.dbg_adr = 32'h23978; force soc.dbg_do = 32'h00c6d533; #1000;
force soc.dbg_adr = 32'h2397c; force soc.dbg_do = 32'h00a7e533; #1000;
force soc.dbg_adr = 32'h23980; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h23984; force soc.dbg_do = 32'h41300693; #1000;
force soc.dbg_adr = 32'h23988; force soc.dbg_do = 32'h40e68733; #1000;
force soc.dbg_adr = 32'h2398c; force soc.dbg_do = 32'h00e7d533; #1000;
force soc.dbg_adr = 32'h23990; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h23994; force soc.dbg_do = 32'h00000513; #1000;
force soc.dbg_adr = 32'h23998; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h2399c; force soc.dbg_do = 32'hfe010113; #1000;
force soc.dbg_adr = 32'h239a0; force soc.dbg_do = 32'h00112e23; #1000;
force soc.dbg_adr = 32'h239a4; force soc.dbg_do = 32'h00812c23; #1000;
force soc.dbg_adr = 32'h239a8; force soc.dbg_do = 32'h00912a23; #1000;
force soc.dbg_adr = 32'h239ac; force soc.dbg_do = 32'h01212823; #1000;
force soc.dbg_adr = 32'h239b0; force soc.dbg_do = 32'h01312623; #1000;
force soc.dbg_adr = 32'h239b4; force soc.dbg_do = 32'h00050793; #1000;
force soc.dbg_adr = 32'h239b8; force soc.dbg_do = 32'h08050663; #1000;
force soc.dbg_adr = 32'h239bc; force soc.dbg_do = 32'h41f55713; #1000;
force soc.dbg_adr = 32'h239c0; force soc.dbg_do = 32'h00a74933; #1000;
force soc.dbg_adr = 32'h239c4; force soc.dbg_do = 32'h40e90933; #1000;
force soc.dbg_adr = 32'h239c8; force soc.dbg_do = 32'h01f55993; #1000;
force soc.dbg_adr = 32'h239cc; force soc.dbg_do = 32'h00090513; #1000;
force soc.dbg_adr = 32'h239d0; force soc.dbg_do = 32'h158000ef; #1000;
force soc.dbg_adr = 32'h239d4; force soc.dbg_do = 32'h41e00793; #1000;
force soc.dbg_adr = 32'h239d8; force soc.dbg_do = 32'h00a00713; #1000;
force soc.dbg_adr = 32'h239dc; force soc.dbg_do = 32'h40a787b3; #1000;
force soc.dbg_adr = 32'h239e0; force soc.dbg_do = 32'h04a74a63; #1000;
force soc.dbg_adr = 32'h239e4; force soc.dbg_do = 32'h00b00713; #1000;
force soc.dbg_adr = 32'h239e8; force soc.dbg_do = 32'h40a70733; #1000;
force soc.dbg_adr = 32'h239ec; force soc.dbg_do = 32'h01550513; #1000;
force soc.dbg_adr = 32'h239f0; force soc.dbg_do = 32'h00e95733; #1000;
force soc.dbg_adr = 32'h239f4; force soc.dbg_do = 32'h00a91933; #1000;
force soc.dbg_adr = 32'h239f8; force soc.dbg_do = 32'h00c71713; #1000;
force soc.dbg_adr = 32'h239fc; force soc.dbg_do = 32'h01c12083; #1000;
force soc.dbg_adr = 32'h23a00; force soc.dbg_do = 32'h01812403; #1000;
force soc.dbg_adr = 32'h23a04; force soc.dbg_do = 32'h00c75713; #1000;
force soc.dbg_adr = 32'h23a08; force soc.dbg_do = 32'h01479793; #1000;
force soc.dbg_adr = 32'h23a0c; force soc.dbg_do = 32'h01f99993; #1000;
force soc.dbg_adr = 32'h23a10; force soc.dbg_do = 32'h00e7e7b3; #1000;
force soc.dbg_adr = 32'h23a14; force soc.dbg_do = 32'h0137e733; #1000;
force soc.dbg_adr = 32'h23a18; force soc.dbg_do = 32'h01412483; #1000;
force soc.dbg_adr = 32'h23a1c; force soc.dbg_do = 32'h00c12983; #1000;
force soc.dbg_adr = 32'h23a20; force soc.dbg_do = 32'h00090513; #1000;
force soc.dbg_adr = 32'h23a24; force soc.dbg_do = 32'h00070593; #1000;
force soc.dbg_adr = 32'h23a28; force soc.dbg_do = 32'h01012903; #1000;
force soc.dbg_adr = 32'h23a2c; force soc.dbg_do = 32'h02010113; #1000;
force soc.dbg_adr = 32'h23a30; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h23a34; force soc.dbg_do = 32'hff550513; #1000;
force soc.dbg_adr = 32'h23a38; force soc.dbg_do = 32'h00a91733; #1000;
force soc.dbg_adr = 32'h23a3c; force soc.dbg_do = 32'h00000913; #1000;
force soc.dbg_adr = 32'h23a40; force soc.dbg_do = 32'hfb9ff06f; #1000;
force soc.dbg_adr = 32'h23a44; force soc.dbg_do = 32'h00000993; #1000;
force soc.dbg_adr = 32'h23a48; force soc.dbg_do = 32'h00000713; #1000;
force soc.dbg_adr = 32'h23a4c; force soc.dbg_do = 32'hff1ff06f; #1000;
force soc.dbg_adr = 32'h23a50; force soc.dbg_do = 32'h00050613; #1000;
force soc.dbg_adr = 32'h23a54; force soc.dbg_do = 32'h00000513; #1000;
force soc.dbg_adr = 32'h23a58; force soc.dbg_do = 32'h0015f693; #1000;
force soc.dbg_adr = 32'h23a5c; force soc.dbg_do = 32'h00068463; #1000;
force soc.dbg_adr = 32'h23a60; force soc.dbg_do = 32'h00c50533; #1000;
force soc.dbg_adr = 32'h23a64; force soc.dbg_do = 32'h0015d593; #1000;
force soc.dbg_adr = 32'h23a68; force soc.dbg_do = 32'h00161613; #1000;
force soc.dbg_adr = 32'h23a6c; force soc.dbg_do = 32'hfe0596e3; #1000;
force soc.dbg_adr = 32'h23a70; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h23a74; force soc.dbg_do = 32'h06054063; #1000;
force soc.dbg_adr = 32'h23a78; force soc.dbg_do = 32'h0605c663; #1000;
force soc.dbg_adr = 32'h23a7c; force soc.dbg_do = 32'h00058613; #1000;
force soc.dbg_adr = 32'h23a80; force soc.dbg_do = 32'h00050593; #1000;
force soc.dbg_adr = 32'h23a84; force soc.dbg_do = 32'hfff00513; #1000;
force soc.dbg_adr = 32'h23a88; force soc.dbg_do = 32'h02060c63; #1000;
force soc.dbg_adr = 32'h23a8c; force soc.dbg_do = 32'h00100693; #1000;
force soc.dbg_adr = 32'h23a90; force soc.dbg_do = 32'h00b67a63; #1000;
force soc.dbg_adr = 32'h23a94; force soc.dbg_do = 32'h00c05863; #1000;
force soc.dbg_adr = 32'h23a98; force soc.dbg_do = 32'h00161613; #1000;
force soc.dbg_adr = 32'h23a9c; force soc.dbg_do = 32'h00169693; #1000;
force soc.dbg_adr = 32'h23aa0; force soc.dbg_do = 32'hfeb66ae3; #1000;
force soc.dbg_adr = 32'h23aa4; force soc.dbg_do = 32'h00000513; #1000;
force soc.dbg_adr = 32'h23aa8; force soc.dbg_do = 32'h00c5e663; #1000;
force soc.dbg_adr = 32'h23aac; force soc.dbg_do = 32'h40c585b3; #1000;
force soc.dbg_adr = 32'h23ab0; force soc.dbg_do = 32'h00d56533; #1000;
force soc.dbg_adr = 32'h23ab4; force soc.dbg_do = 32'h0016d693; #1000;
force soc.dbg_adr = 32'h23ab8; force soc.dbg_do = 32'h00165613; #1000;
force soc.dbg_adr = 32'h23abc; force soc.dbg_do = 32'hfe0696e3; #1000;
force soc.dbg_adr = 32'h23ac0; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h23ac4; force soc.dbg_do = 32'h00008293; #1000;
force soc.dbg_adr = 32'h23ac8; force soc.dbg_do = 32'hfb5ff0ef; #1000;
force soc.dbg_adr = 32'h23acc; force soc.dbg_do = 32'h00058513; #1000;
force soc.dbg_adr = 32'h23ad0; force soc.dbg_do = 32'h00028067; #1000;
force soc.dbg_adr = 32'h23ad4; force soc.dbg_do = 32'h40a00533; #1000;
force soc.dbg_adr = 32'h23ad8; force soc.dbg_do = 32'h00b04863; #1000;
force soc.dbg_adr = 32'h23adc; force soc.dbg_do = 32'h40b005b3; #1000;
force soc.dbg_adr = 32'h23ae0; force soc.dbg_do = 32'hf9dff06f; #1000;
force soc.dbg_adr = 32'h23ae4; force soc.dbg_do = 32'h40b005b3; #1000;
force soc.dbg_adr = 32'h23ae8; force soc.dbg_do = 32'h00008293; #1000;
force soc.dbg_adr = 32'h23aec; force soc.dbg_do = 32'hf91ff0ef; #1000;
force soc.dbg_adr = 32'h23af0; force soc.dbg_do = 32'h40a00533; #1000;
force soc.dbg_adr = 32'h23af4; force soc.dbg_do = 32'h00028067; #1000;
force soc.dbg_adr = 32'h23af8; force soc.dbg_do = 32'h00008293; #1000;
force soc.dbg_adr = 32'h23afc; force soc.dbg_do = 32'h0005ca63; #1000;
force soc.dbg_adr = 32'h23b00; force soc.dbg_do = 32'h00054c63; #1000;
force soc.dbg_adr = 32'h23b04; force soc.dbg_do = 32'hf79ff0ef; #1000;
force soc.dbg_adr = 32'h23b08; force soc.dbg_do = 32'h00058513; #1000;
force soc.dbg_adr = 32'h23b0c; force soc.dbg_do = 32'h00028067; #1000;
force soc.dbg_adr = 32'h23b10; force soc.dbg_do = 32'h40b005b3; #1000;
force soc.dbg_adr = 32'h23b14; force soc.dbg_do = 32'hfe0558e3; #1000;
force soc.dbg_adr = 32'h23b18; force soc.dbg_do = 32'h40a00533; #1000;
force soc.dbg_adr = 32'h23b1c; force soc.dbg_do = 32'hf61ff0ef; #1000;
force soc.dbg_adr = 32'h23b20; force soc.dbg_do = 32'h40b00533; #1000;
force soc.dbg_adr = 32'h23b24; force soc.dbg_do = 32'h00028067; #1000;
force soc.dbg_adr = 32'h23b28; force soc.dbg_do = 32'h000107b7; #1000;
force soc.dbg_adr = 32'h23b2c; force soc.dbg_do = 32'h02f57a63; #1000;
force soc.dbg_adr = 32'h23b30; force soc.dbg_do = 32'h10053793; #1000;
force soc.dbg_adr = 32'h23b34; force soc.dbg_do = 32'h0017b793; #1000;
force soc.dbg_adr = 32'h23b38; force soc.dbg_do = 32'h00379793; #1000;
force soc.dbg_adr = 32'h23b3c; force soc.dbg_do = 32'h00024737; #1000;
force soc.dbg_adr = 32'h23b40; force soc.dbg_do = 32'h02000693; #1000;
force soc.dbg_adr = 32'h23b44; force soc.dbg_do = 32'h40f686b3; #1000;
force soc.dbg_adr = 32'h23b48; force soc.dbg_do = 32'h00f55533; #1000;
force soc.dbg_adr = 32'h23b4c; force soc.dbg_do = 32'h20870793; #1000;
force soc.dbg_adr = 32'h23b50; force soc.dbg_do = 32'h00a787b3; #1000;
force soc.dbg_adr = 32'h23b54; force soc.dbg_do = 32'h0007c503; #1000;
force soc.dbg_adr = 32'h23b58; force soc.dbg_do = 32'h40a68533; #1000;
force soc.dbg_adr = 32'h23b5c; force soc.dbg_do = 32'h00008067; #1000;
force soc.dbg_adr = 32'h23b60; force soc.dbg_do = 32'h01000737; #1000;
force soc.dbg_adr = 32'h23b64; force soc.dbg_do = 32'h01800793; #1000;
force soc.dbg_adr = 32'h23b68; force soc.dbg_do = 32'hfce57ae3; #1000;
force soc.dbg_adr = 32'h23b6c; force soc.dbg_do = 32'h01000793; #1000;
force soc.dbg_adr = 32'h23b70; force soc.dbg_do = 32'hfcdff06f; #1000;
force soc.dbg_adr = 32'h23b74; force soc.dbg_do = 32'h20737362; #1000;
force soc.dbg_adr = 32'h23b78; force soc.dbg_do = 32'h203a7025; #1000;
force soc.dbg_adr = 32'h23b7c; force soc.dbg_do = 32'h000a6425; #1000;
force soc.dbg_adr = 32'h23b80; force soc.dbg_do = 32'h736e7572; #1000;
force soc.dbg_adr = 32'h23b84; force soc.dbg_do = 32'h2020203a; #1000;
force soc.dbg_adr = 32'h23b88; force soc.dbg_do = 32'h000a6425; #1000;
force soc.dbg_adr = 32'h23b8c; force soc.dbg_do = 32'h6c637963; #1000;
force soc.dbg_adr = 32'h23b90; force soc.dbg_do = 32'h203a7365; #1000;
force soc.dbg_adr = 32'h23b94; force soc.dbg_do = 32'h000a6425; #1000;
force soc.dbg_adr = 32'h23b98; force soc.dbg_do = 32'h74736e69; #1000;
force soc.dbg_adr = 32'h23b9c; force soc.dbg_do = 32'h20203a72; #1000;
force soc.dbg_adr = 32'h23ba0; force soc.dbg_do = 32'h000a6425; #1000;
force soc.dbg_adr = 32'h23ba4; force soc.dbg_do = 32'h656d6974; #1000;
force soc.dbg_adr = 32'h23ba8; force soc.dbg_do = 32'h2020203a; #1000;
force soc.dbg_adr = 32'h23bac; force soc.dbg_do = 32'h75206425; #1000;
force soc.dbg_adr = 32'h23bb0; force soc.dbg_do = 32'h25282073; #1000;
force soc.dbg_adr = 32'h23bb4; force soc.dbg_do = 32'h30252e64; #1000;
force soc.dbg_adr = 32'h23bb8; force soc.dbg_do = 32'h73206436; #1000;
force soc.dbg_adr = 32'h23bbc; force soc.dbg_do = 32'h00000a29; #1000;
force soc.dbg_adr = 32'h23bc0; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h23bc4; force soc.dbg_do = 32'h0000000a; #1000;
force soc.dbg_adr = 32'h23bc8; force soc.dbg_do = 32'h3a697063; #1000;
force soc.dbg_adr = 32'h23bcc; force soc.dbg_do = 32'h6c6c2520; #1000;
force soc.dbg_adr = 32'h23bd0; force soc.dbg_do = 32'h30252e75; #1000;
force soc.dbg_adr = 32'h23bd4; force soc.dbg_do = 32'h756c6c33; #1000;
force soc.dbg_adr = 32'h23bd8; force soc.dbg_do = 32'h0000000a; #1000;
force soc.dbg_adr = 32'h23bdc; force soc.dbg_do = 32'h3a637069; #1000;
force soc.dbg_adr = 32'h23be0; force soc.dbg_do = 32'h6c6c2520; #1000;
force soc.dbg_adr = 32'h23be4; force soc.dbg_do = 32'h30252e75; #1000;
force soc.dbg_adr = 32'h23be8; force soc.dbg_do = 32'h756c6c33; #1000;
force soc.dbg_adr = 32'h23bec; force soc.dbg_do = 32'h0000000a; #1000;
force soc.dbg_adr = 32'h23bf0; force soc.dbg_do = 32'h79726864; #1000;
force soc.dbg_adr = 32'h23bf4; force soc.dbg_do = 32'h6e6f7473; #1000;
force soc.dbg_adr = 32'h23bf8; force soc.dbg_do = 32'h70207365; #1000;
force soc.dbg_adr = 32'h23bfc; force soc.dbg_do = 32'h73207265; #1000;
force soc.dbg_adr = 32'h23c00; force soc.dbg_do = 32'h6e6f6365; #1000;
force soc.dbg_adr = 32'h23c04; force soc.dbg_do = 32'h25203a64; #1000;
force soc.dbg_adr = 32'h23c08; force soc.dbg_do = 32'h00000a75; #1000;
force soc.dbg_adr = 32'h23c0c; force soc.dbg_do = 32'h70696d64; #1000;
force soc.dbg_adr = 32'h23c10; force soc.dbg_do = 32'h25203a73; #1000;
force soc.dbg_adr = 32'h23c14; force soc.dbg_do = 32'h30252e64; #1000;
force soc.dbg_adr = 32'h23c18; force soc.dbg_do = 32'h000a6433; #1000;
force soc.dbg_adr = 32'h23c1c; force soc.dbg_do = 32'h70696d64; #1000;
force soc.dbg_adr = 32'h23c20; force soc.dbg_do = 32'h202f2073; #1000;
force soc.dbg_adr = 32'h23c24; force soc.dbg_do = 32'h3a7a484d; #1000;
force soc.dbg_adr = 32'h23c28; force soc.dbg_do = 32'h2e642520; #1000;
force soc.dbg_adr = 32'h23c2c; force soc.dbg_do = 32'h64333025; #1000;
force soc.dbg_adr = 32'h23c30; force soc.dbg_do = 32'h25282020; #1000;
force soc.dbg_adr = 32'h23c34; force soc.dbg_do = 32'h484d2064; #1000;
force soc.dbg_adr = 32'h23c38; force soc.dbg_do = 32'h000a297a; #1000;
force soc.dbg_adr = 32'h23c3c; force soc.dbg_do = 32'h59524844; #1000;
force soc.dbg_adr = 32'h23c40; force soc.dbg_do = 32'h4e4f5453; #1000;
force soc.dbg_adr = 32'h23c44; force soc.dbg_do = 32'h52502045; #1000;
force soc.dbg_adr = 32'h23c48; force soc.dbg_do = 32'h4152474f; #1000;
force soc.dbg_adr = 32'h23c4c; force soc.dbg_do = 32'h53202c4d; #1000;
force soc.dbg_adr = 32'h23c50; force soc.dbg_do = 32'h20454d4f; #1000;
force soc.dbg_adr = 32'h23c54; force soc.dbg_do = 32'h49525453; #1000;
force soc.dbg_adr = 32'h23c58; force soc.dbg_do = 32'h0000474e; #1000;
force soc.dbg_adr = 32'h23c5c; force soc.dbg_do = 32'h59524844; #1000;
force soc.dbg_adr = 32'h23c60; force soc.dbg_do = 32'h4e4f5453; #1000;
force soc.dbg_adr = 32'h23c64; force soc.dbg_do = 32'h52502045; #1000;
force soc.dbg_adr = 32'h23c68; force soc.dbg_do = 32'h4152474f; #1000;
force soc.dbg_adr = 32'h23c6c; force soc.dbg_do = 32'h31202c4d; #1000;
force soc.dbg_adr = 32'h23c70; force soc.dbg_do = 32'h20545327; #1000;
force soc.dbg_adr = 32'h23c74; force soc.dbg_do = 32'h49525453; #1000;
force soc.dbg_adr = 32'h23c78; force soc.dbg_do = 32'h0000474e; #1000;
force soc.dbg_adr = 32'h23c7c; force soc.dbg_do = 32'h79726844; #1000;
force soc.dbg_adr = 32'h23c80; force soc.dbg_do = 32'h6e6f7473; #1000;
force soc.dbg_adr = 32'h23c84; force soc.dbg_do = 32'h65422065; #1000;
force soc.dbg_adr = 32'h23c88; force soc.dbg_do = 32'h6d68636e; #1000;
force soc.dbg_adr = 32'h23c8c; force soc.dbg_do = 32'h2c6b7261; #1000;
force soc.dbg_adr = 32'h23c90; force soc.dbg_do = 32'h72655620; #1000;
force soc.dbg_adr = 32'h23c94; force soc.dbg_do = 32'h6e6f6973; #1000;
force soc.dbg_adr = 32'h23c98; force soc.dbg_do = 32'h312e3220; #1000;
force soc.dbg_adr = 32'h23c9c; force soc.dbg_do = 32'h614c2820; #1000;
force soc.dbg_adr = 32'h23ca0; force soc.dbg_do = 32'h6175676e; #1000;
force soc.dbg_adr = 32'h23ca4; force soc.dbg_do = 32'h203a6567; #1000;
force soc.dbg_adr = 32'h23ca8; force soc.dbg_do = 32'h000a2943; #1000;
force soc.dbg_adr = 32'h23cac; force soc.dbg_do = 32'h676f7250; #1000;
force soc.dbg_adr = 32'h23cb0; force soc.dbg_do = 32'h206d6172; #1000;
force soc.dbg_adr = 32'h23cb4; force soc.dbg_do = 32'h706d6f63; #1000;
force soc.dbg_adr = 32'h23cb8; force soc.dbg_do = 32'h64656c69; #1000;
force soc.dbg_adr = 32'h23cbc; force soc.dbg_do = 32'h74697720; #1000;
force soc.dbg_adr = 32'h23cc0; force soc.dbg_do = 32'h72272068; #1000;
force soc.dbg_adr = 32'h23cc4; force soc.dbg_do = 32'h73696765; #1000;
force soc.dbg_adr = 32'h23cc8; force soc.dbg_do = 32'h27726574; #1000;
force soc.dbg_adr = 32'h23ccc; force soc.dbg_do = 32'h74746120; #1000;
force soc.dbg_adr = 32'h23cd0; force soc.dbg_do = 32'h75626972; #1000;
force soc.dbg_adr = 32'h23cd4; force soc.dbg_do = 32'h000a6574; #1000;
force soc.dbg_adr = 32'h23cd8; force soc.dbg_do = 32'h676f7250; #1000;
force soc.dbg_adr = 32'h23cdc; force soc.dbg_do = 32'h206d6172; #1000;
force soc.dbg_adr = 32'h23ce0; force soc.dbg_do = 32'h706d6f63; #1000;
force soc.dbg_adr = 32'h23ce4; force soc.dbg_do = 32'h64656c69; #1000;
force soc.dbg_adr = 32'h23ce8; force soc.dbg_do = 32'h74697720; #1000;
force soc.dbg_adr = 32'h23cec; force soc.dbg_do = 32'h74756f68; #1000;
force soc.dbg_adr = 32'h23cf0; force soc.dbg_do = 32'h65722720; #1000;
force soc.dbg_adr = 32'h23cf4; force soc.dbg_do = 32'h74736967; #1000;
force soc.dbg_adr = 32'h23cf8; force soc.dbg_do = 32'h20277265; #1000;
force soc.dbg_adr = 32'h23cfc; force soc.dbg_do = 32'h72747461; #1000;
force soc.dbg_adr = 32'h23d00; force soc.dbg_do = 32'h74756269; #1000;
force soc.dbg_adr = 32'h23d04; force soc.dbg_do = 32'h00000a65; #1000;
force soc.dbg_adr = 32'h23d08; force soc.dbg_do = 32'h63657845; #1000;
force soc.dbg_adr = 32'h23d0c; force soc.dbg_do = 32'h6f697475; #1000;
force soc.dbg_adr = 32'h23d10; force soc.dbg_do = 32'h7473206e; #1000;
force soc.dbg_adr = 32'h23d14; force soc.dbg_do = 32'h73747261; #1000;
force soc.dbg_adr = 32'h23d18; force soc.dbg_do = 32'h6425202c; #1000;
force soc.dbg_adr = 32'h23d1c; force soc.dbg_do = 32'h6e757220; #1000;
force soc.dbg_adr = 32'h23d20; force soc.dbg_do = 32'h68742073; #1000;
force soc.dbg_adr = 32'h23d24; force soc.dbg_do = 32'h67756f72; #1000;
force soc.dbg_adr = 32'h23d28; force soc.dbg_do = 32'h68442068; #1000;
force soc.dbg_adr = 32'h23d2c; force soc.dbg_do = 32'h74737972; #1000;
force soc.dbg_adr = 32'h23d30; force soc.dbg_do = 32'h0a656e6f; #1000;
force soc.dbg_adr = 32'h23d34; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h23d38; force soc.dbg_do = 32'h59524844; #1000;
force soc.dbg_adr = 32'h23d3c; force soc.dbg_do = 32'h4e4f5453; #1000;
force soc.dbg_adr = 32'h23d40; force soc.dbg_do = 32'h52502045; #1000;
force soc.dbg_adr = 32'h23d44; force soc.dbg_do = 32'h4152474f; #1000;
force soc.dbg_adr = 32'h23d48; force soc.dbg_do = 32'h32202c4d; #1000;
force soc.dbg_adr = 32'h23d4c; force soc.dbg_do = 32'h20444e27; #1000;
force soc.dbg_adr = 32'h23d50; force soc.dbg_do = 32'h49525453; #1000;
force soc.dbg_adr = 32'h23d54; force soc.dbg_do = 32'h0000474e; #1000;
force soc.dbg_adr = 32'h23d58; force soc.dbg_do = 32'h59524844; #1000;
force soc.dbg_adr = 32'h23d5c; force soc.dbg_do = 32'h4e4f5453; #1000;
force soc.dbg_adr = 32'h23d60; force soc.dbg_do = 32'h52502045; #1000;
force soc.dbg_adr = 32'h23d64; force soc.dbg_do = 32'h4152474f; #1000;
force soc.dbg_adr = 32'h23d68; force soc.dbg_do = 32'h33202c4d; #1000;
force soc.dbg_adr = 32'h23d6c; force soc.dbg_do = 32'h20445227; #1000;
force soc.dbg_adr = 32'h23d70; force soc.dbg_do = 32'h49525453; #1000;
force soc.dbg_adr = 32'h23d74; force soc.dbg_do = 32'h0000474e; #1000;
force soc.dbg_adr = 32'h23d78; force soc.dbg_do = 32'h63657845; #1000;
force soc.dbg_adr = 32'h23d7c; force soc.dbg_do = 32'h6f697475; #1000;
force soc.dbg_adr = 32'h23d80; force soc.dbg_do = 32'h6e65206e; #1000;
force soc.dbg_adr = 32'h23d84; force soc.dbg_do = 32'h000a7364; #1000;
force soc.dbg_adr = 32'h23d88; force soc.dbg_do = 32'h616e6946; #1000;
force soc.dbg_adr = 32'h23d8c; force soc.dbg_do = 32'h6176206c; #1000;
force soc.dbg_adr = 32'h23d90; force soc.dbg_do = 32'h7365756c; #1000;
force soc.dbg_adr = 32'h23d94; force soc.dbg_do = 32'h20666f20; #1000;
force soc.dbg_adr = 32'h23d98; force soc.dbg_do = 32'h20656874; #1000;
force soc.dbg_adr = 32'h23d9c; force soc.dbg_do = 32'h69726176; #1000;
force soc.dbg_adr = 32'h23da0; force soc.dbg_do = 32'h656c6261; #1000;
force soc.dbg_adr = 32'h23da4; force soc.dbg_do = 32'h73752073; #1000;
force soc.dbg_adr = 32'h23da8; force soc.dbg_do = 32'h69206465; #1000;
force soc.dbg_adr = 32'h23dac; force soc.dbg_do = 32'h6874206e; #1000;
force soc.dbg_adr = 32'h23db0; force soc.dbg_do = 32'h65622065; #1000;
force soc.dbg_adr = 32'h23db4; force soc.dbg_do = 32'h6d68636e; #1000;
force soc.dbg_adr = 32'h23db8; force soc.dbg_do = 32'h3a6b7261; #1000;
force soc.dbg_adr = 32'h23dbc; force soc.dbg_do = 32'h0000000a; #1000;
force soc.dbg_adr = 32'h23dc0; force soc.dbg_do = 32'h5f746e49; #1000;
force soc.dbg_adr = 32'h23dc4; force soc.dbg_do = 32'h626f6c47; #1000;
force soc.dbg_adr = 32'h23dc8; force soc.dbg_do = 32'h2020203a; #1000;
force soc.dbg_adr = 32'h23dcc; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23dd0; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23dd4; force soc.dbg_do = 32'h0a642520; #1000;
force soc.dbg_adr = 32'h23dd8; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h23ddc; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23de0; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23de4; force soc.dbg_do = 32'h756f6873; #1000;
force soc.dbg_adr = 32'h23de8; force soc.dbg_do = 32'h6220646c; #1000;
force soc.dbg_adr = 32'h23dec; force soc.dbg_do = 32'h20203a65; #1000;
force soc.dbg_adr = 32'h23df0; force soc.dbg_do = 32'h0a642520; #1000;
force soc.dbg_adr = 32'h23df4; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h23df8; force soc.dbg_do = 32'h6c6f6f42; #1000;
force soc.dbg_adr = 32'h23dfc; force soc.dbg_do = 32'h6f6c475f; #1000;
force soc.dbg_adr = 32'h23e00; force soc.dbg_do = 32'h20203a62; #1000;
force soc.dbg_adr = 32'h23e04; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23e08; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23e0c; force soc.dbg_do = 32'h0a642520; #1000;
force soc.dbg_adr = 32'h23e10; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h23e14; force soc.dbg_do = 32'h315f6843; #1000;
force soc.dbg_adr = 32'h23e18; force soc.dbg_do = 32'h6f6c475f; #1000;
force soc.dbg_adr = 32'h23e1c; force soc.dbg_do = 32'h20203a62; #1000;
force soc.dbg_adr = 32'h23e20; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23e24; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23e28; force soc.dbg_do = 32'h0a632520; #1000;
force soc.dbg_adr = 32'h23e2c; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h23e30; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23e34; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23e38; force soc.dbg_do = 32'h756f6873; #1000;
force soc.dbg_adr = 32'h23e3c; force soc.dbg_do = 32'h6220646c; #1000;
force soc.dbg_adr = 32'h23e40; force soc.dbg_do = 32'h20203a65; #1000;
force soc.dbg_adr = 32'h23e44; force soc.dbg_do = 32'h0a632520; #1000;
force soc.dbg_adr = 32'h23e48; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h23e4c; force soc.dbg_do = 32'h325f6843; #1000;
force soc.dbg_adr = 32'h23e50; force soc.dbg_do = 32'h6f6c475f; #1000;
force soc.dbg_adr = 32'h23e54; force soc.dbg_do = 32'h20203a62; #1000;
force soc.dbg_adr = 32'h23e58; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23e5c; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23e60; force soc.dbg_do = 32'h0a632520; #1000;
force soc.dbg_adr = 32'h23e64; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h23e68; force soc.dbg_do = 32'h5f727241; #1000;
force soc.dbg_adr = 32'h23e6c; force soc.dbg_do = 32'h6c475f31; #1000;
force soc.dbg_adr = 32'h23e70; force soc.dbg_do = 32'h385b626f; #1000;
force soc.dbg_adr = 32'h23e74; force soc.dbg_do = 32'h20203a5d; #1000;
force soc.dbg_adr = 32'h23e78; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23e7c; force soc.dbg_do = 32'h0a642520; #1000;
force soc.dbg_adr = 32'h23e80; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h23e84; force soc.dbg_do = 32'h5f727241; #1000;
force soc.dbg_adr = 32'h23e88; force soc.dbg_do = 32'h6c475f32; #1000;
force soc.dbg_adr = 32'h23e8c; force soc.dbg_do = 32'h385b626f; #1000;
force soc.dbg_adr = 32'h23e90; force soc.dbg_do = 32'h5d375b5d; #1000;
force soc.dbg_adr = 32'h23e94; force soc.dbg_do = 32'h2020203a; #1000;
force soc.dbg_adr = 32'h23e98; force soc.dbg_do = 32'h0a642520; #1000;
force soc.dbg_adr = 32'h23e9c; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h23ea0; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23ea4; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23ea8; force soc.dbg_do = 32'h756f6873; #1000;
force soc.dbg_adr = 32'h23eac; force soc.dbg_do = 32'h6220646c; #1000;
force soc.dbg_adr = 32'h23eb0; force soc.dbg_do = 32'h20203a65; #1000;
force soc.dbg_adr = 32'h23eb4; force soc.dbg_do = 32'h6d754e20; #1000;
force soc.dbg_adr = 32'h23eb8; force soc.dbg_do = 32'h5f726562; #1000;
force soc.dbg_adr = 32'h23ebc; force soc.dbg_do = 32'h525f664f; #1000;
force soc.dbg_adr = 32'h23ec0; force soc.dbg_do = 32'h20736e75; #1000;
force soc.dbg_adr = 32'h23ec4; force soc.dbg_do = 32'h3031202b; #1000;
force soc.dbg_adr = 32'h23ec8; force soc.dbg_do = 32'h0000000a; #1000;
force soc.dbg_adr = 32'h23ecc; force soc.dbg_do = 32'h5f727450; #1000;
force soc.dbg_adr = 32'h23ed0; force soc.dbg_do = 32'h626f6c47; #1000;
force soc.dbg_adr = 32'h23ed4; force soc.dbg_do = 32'h000a3e2d; #1000;
force soc.dbg_adr = 32'h23ed8; force soc.dbg_do = 32'h74502020; #1000;
force soc.dbg_adr = 32'h23edc; force soc.dbg_do = 32'h6f435f72; #1000;
force soc.dbg_adr = 32'h23ee0; force soc.dbg_do = 32'h203a706d; #1000;
force soc.dbg_adr = 32'h23ee4; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23ee8; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23eec; force soc.dbg_do = 32'h0a642520; #1000;
force soc.dbg_adr = 32'h23ef0; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h23ef4; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23ef8; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23efc; force soc.dbg_do = 32'h756f6873; #1000;
force soc.dbg_adr = 32'h23f00; force soc.dbg_do = 32'h6220646c; #1000;
force soc.dbg_adr = 32'h23f04; force soc.dbg_do = 32'h20203a65; #1000;
force soc.dbg_adr = 32'h23f08; force soc.dbg_do = 32'h6d692820; #1000;
force soc.dbg_adr = 32'h23f0c; force soc.dbg_do = 32'h6d656c70; #1000;
force soc.dbg_adr = 32'h23f10; force soc.dbg_do = 32'h61746e65; #1000;
force soc.dbg_adr = 32'h23f14; force soc.dbg_do = 32'h6e6f6974; #1000;
force soc.dbg_adr = 32'h23f18; force soc.dbg_do = 32'h7065642d; #1000;
force soc.dbg_adr = 32'h23f1c; force soc.dbg_do = 32'h65646e65; #1000;
force soc.dbg_adr = 32'h23f20; force soc.dbg_do = 32'h0a29746e; #1000;
force soc.dbg_adr = 32'h23f24; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h23f28; force soc.dbg_do = 32'h69442020; #1000;
force soc.dbg_adr = 32'h23f2c; force soc.dbg_do = 32'h3a726373; #1000;
force soc.dbg_adr = 32'h23f30; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23f34; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23f38; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23f3c; force soc.dbg_do = 32'h0a642520; #1000;
force soc.dbg_adr = 32'h23f40; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h23f44; force soc.dbg_do = 32'h6e452020; #1000;
force soc.dbg_adr = 32'h23f48; force soc.dbg_do = 32'h435f6d75; #1000;
force soc.dbg_adr = 32'h23f4c; force soc.dbg_do = 32'h3a706d6f; #1000;
force soc.dbg_adr = 32'h23f50; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23f54; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23f58; force soc.dbg_do = 32'h0a642520; #1000;
force soc.dbg_adr = 32'h23f5c; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h23f60; force soc.dbg_do = 32'h6e492020; #1000;
force soc.dbg_adr = 32'h23f64; force soc.dbg_do = 32'h6f435f74; #1000;
force soc.dbg_adr = 32'h23f68; force soc.dbg_do = 32'h203a706d; #1000;
force soc.dbg_adr = 32'h23f6c; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23f70; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23f74; force soc.dbg_do = 32'h0a642520; #1000;
force soc.dbg_adr = 32'h23f78; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h23f7c; force soc.dbg_do = 32'h74532020; #1000;
force soc.dbg_adr = 32'h23f80; force soc.dbg_do = 32'h6f435f72; #1000;
force soc.dbg_adr = 32'h23f84; force soc.dbg_do = 32'h203a706d; #1000;
force soc.dbg_adr = 32'h23f88; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23f8c; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23f90; force soc.dbg_do = 32'h0a732520; #1000;
force soc.dbg_adr = 32'h23f94; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h23f98; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23f9c; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23fa0; force soc.dbg_do = 32'h756f6873; #1000;
force soc.dbg_adr = 32'h23fa4; force soc.dbg_do = 32'h6220646c; #1000;
force soc.dbg_adr = 32'h23fa8; force soc.dbg_do = 32'h20203a65; #1000;
force soc.dbg_adr = 32'h23fac; force soc.dbg_do = 32'h52484420; #1000;
force soc.dbg_adr = 32'h23fb0; force soc.dbg_do = 32'h4f545359; #1000;
force soc.dbg_adr = 32'h23fb4; force soc.dbg_do = 32'h5020454e; #1000;
force soc.dbg_adr = 32'h23fb8; force soc.dbg_do = 32'h52474f52; #1000;
force soc.dbg_adr = 32'h23fbc; force soc.dbg_do = 32'h202c4d41; #1000;
force soc.dbg_adr = 32'h23fc0; force soc.dbg_do = 32'h454d4f53; #1000;
force soc.dbg_adr = 32'h23fc4; force soc.dbg_do = 32'h52545320; #1000;
force soc.dbg_adr = 32'h23fc8; force soc.dbg_do = 32'h0a474e49; #1000;
force soc.dbg_adr = 32'h23fcc; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h23fd0; force soc.dbg_do = 32'h7478654e; #1000;
force soc.dbg_adr = 32'h23fd4; force soc.dbg_do = 32'h7274505f; #1000;
force soc.dbg_adr = 32'h23fd8; force soc.dbg_do = 32'h6f6c475f; #1000;
force soc.dbg_adr = 32'h23fdc; force soc.dbg_do = 32'h0a3e2d62; #1000;
force soc.dbg_adr = 32'h23fe0; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h23fe4; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23fe8; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h23fec; force soc.dbg_do = 32'h756f6873; #1000;
force soc.dbg_adr = 32'h23ff0; force soc.dbg_do = 32'h6220646c; #1000;
force soc.dbg_adr = 32'h23ff4; force soc.dbg_do = 32'h20203a65; #1000;
force soc.dbg_adr = 32'h23ff8; force soc.dbg_do = 32'h6d692820; #1000;
force soc.dbg_adr = 32'h23ffc; force soc.dbg_do = 32'h6d656c70; #1000;
force soc.dbg_adr = 32'h24000; force soc.dbg_do = 32'h61746e65; #1000;
force soc.dbg_adr = 32'h24004; force soc.dbg_do = 32'h6e6f6974; #1000;
force soc.dbg_adr = 32'h24008; force soc.dbg_do = 32'h7065642d; #1000;
force soc.dbg_adr = 32'h2400c; force soc.dbg_do = 32'h65646e65; #1000;
force soc.dbg_adr = 32'h24010; force soc.dbg_do = 32'h2c29746e; #1000;
force soc.dbg_adr = 32'h24014; force soc.dbg_do = 32'h6d617320; #1000;
force soc.dbg_adr = 32'h24018; force soc.dbg_do = 32'h73612065; #1000;
force soc.dbg_adr = 32'h2401c; force soc.dbg_do = 32'h6f626120; #1000;
force soc.dbg_adr = 32'h24020; force soc.dbg_do = 32'h000a6576; #1000;
force soc.dbg_adr = 32'h24024; force soc.dbg_do = 32'h5f746e49; #1000;
force soc.dbg_adr = 32'h24028; force soc.dbg_do = 32'h6f4c5f31; #1000;
force soc.dbg_adr = 32'h2402c; force soc.dbg_do = 32'h20203a63; #1000;
force soc.dbg_adr = 32'h24030; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h24034; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h24038; force soc.dbg_do = 32'h0a642520; #1000;
force soc.dbg_adr = 32'h2403c; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h24040; force soc.dbg_do = 32'h5f746e49; #1000;
force soc.dbg_adr = 32'h24044; force soc.dbg_do = 32'h6f4c5f32; #1000;
force soc.dbg_adr = 32'h24048; force soc.dbg_do = 32'h20203a63; #1000;
force soc.dbg_adr = 32'h2404c; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h24050; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h24054; force soc.dbg_do = 32'h0a642520; #1000;
force soc.dbg_adr = 32'h24058; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h2405c; force soc.dbg_do = 32'h5f746e49; #1000;
force soc.dbg_adr = 32'h24060; force soc.dbg_do = 32'h6f4c5f33; #1000;
force soc.dbg_adr = 32'h24064; force soc.dbg_do = 32'h20203a63; #1000;
force soc.dbg_adr = 32'h24068; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h2406c; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h24070; force soc.dbg_do = 32'h0a642520; #1000;
force soc.dbg_adr = 32'h24074; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h24078; force soc.dbg_do = 32'h6d756e45; #1000;
force soc.dbg_adr = 32'h2407c; force soc.dbg_do = 32'h636f4c5f; #1000;
force soc.dbg_adr = 32'h24080; force soc.dbg_do = 32'h2020203a; #1000;
force soc.dbg_adr = 32'h24084; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h24088; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h2408c; force soc.dbg_do = 32'h0a642520; #1000;
force soc.dbg_adr = 32'h24090; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h24094; force soc.dbg_do = 32'h5f727453; #1000;
force soc.dbg_adr = 32'h24098; force soc.dbg_do = 32'h6f4c5f31; #1000;
force soc.dbg_adr = 32'h2409c; force soc.dbg_do = 32'h20203a63; #1000;
force soc.dbg_adr = 32'h240a0; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h240a4; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h240a8; force soc.dbg_do = 32'h0a732520; #1000;
force soc.dbg_adr = 32'h240ac; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h240b0; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h240b4; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h240b8; force soc.dbg_do = 32'h756f6873; #1000;
force soc.dbg_adr = 32'h240bc; force soc.dbg_do = 32'h6220646c; #1000;
force soc.dbg_adr = 32'h240c0; force soc.dbg_do = 32'h20203a65; #1000;
force soc.dbg_adr = 32'h240c4; force soc.dbg_do = 32'h52484420; #1000;
force soc.dbg_adr = 32'h240c8; force soc.dbg_do = 32'h4f545359; #1000;
force soc.dbg_adr = 32'h240cc; force soc.dbg_do = 32'h5020454e; #1000;
force soc.dbg_adr = 32'h240d0; force soc.dbg_do = 32'h52474f52; #1000;
force soc.dbg_adr = 32'h240d4; force soc.dbg_do = 32'h202c4d41; #1000;
force soc.dbg_adr = 32'h240d8; force soc.dbg_do = 32'h54532731; #1000;
force soc.dbg_adr = 32'h240dc; force soc.dbg_do = 32'h52545320; #1000;
force soc.dbg_adr = 32'h240e0; force soc.dbg_do = 32'h0a474e49; #1000;
force soc.dbg_adr = 32'h240e4; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h240e8; force soc.dbg_do = 32'h5f727453; #1000;
force soc.dbg_adr = 32'h240ec; force soc.dbg_do = 32'h6f4c5f32; #1000;
force soc.dbg_adr = 32'h240f0; force soc.dbg_do = 32'h20203a63; #1000;
force soc.dbg_adr = 32'h240f4; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h240f8; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h240fc; force soc.dbg_do = 32'h0a732520; #1000;
force soc.dbg_adr = 32'h24100; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h24104; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h24108; force soc.dbg_do = 32'h20202020; #1000;
force soc.dbg_adr = 32'h2410c; force soc.dbg_do = 32'h756f6873; #1000;
force soc.dbg_adr = 32'h24110; force soc.dbg_do = 32'h6220646c; #1000;
force soc.dbg_adr = 32'h24114; force soc.dbg_do = 32'h20203a65; #1000;
force soc.dbg_adr = 32'h24118; force soc.dbg_do = 32'h52484420; #1000;
force soc.dbg_adr = 32'h2411c; force soc.dbg_do = 32'h4f545359; #1000;
force soc.dbg_adr = 32'h24120; force soc.dbg_do = 32'h5020454e; #1000;
force soc.dbg_adr = 32'h24124; force soc.dbg_do = 32'h52474f52; #1000;
force soc.dbg_adr = 32'h24128; force soc.dbg_do = 32'h202c4d41; #1000;
force soc.dbg_adr = 32'h2412c; force soc.dbg_do = 32'h444e2732; #1000;
force soc.dbg_adr = 32'h24130; force soc.dbg_do = 32'h52545320; #1000;
force soc.dbg_adr = 32'h24134; force soc.dbg_do = 32'h0a474e49; #1000;
force soc.dbg_adr = 32'h24138; force soc.dbg_do = 32'h00000000; #1000;
force soc.dbg_adr = 32'h2413c; force soc.dbg_do = 32'h00021720; #1000;
force soc.dbg_adr = 32'h24140; force soc.dbg_do = 32'h000216a4; #1000;
force soc.dbg_adr = 32'h24144; force soc.dbg_do = 32'h000216a4; #1000;
force soc.dbg_adr = 32'h24148; force soc.dbg_do = 32'h00021714; #1000;
force soc.dbg_adr = 32'h2414c; force soc.dbg_do = 32'h000216a4; #1000;
force soc.dbg_adr = 32'h24150; force soc.dbg_do = 32'h000216a4; #1000;
force soc.dbg_adr = 32'h24154; force soc.dbg_do = 32'h000216a4; #1000;
force soc.dbg_adr = 32'h24158; force soc.dbg_do = 32'h000216a4; #1000;
force soc.dbg_adr = 32'h2415c; force soc.dbg_do = 32'h000216a4; #1000;
force soc.dbg_adr = 32'h24160; force soc.dbg_do = 32'h000216a4; #1000;
force soc.dbg_adr = 32'h24164; force soc.dbg_do = 32'h000216a4; #1000;
force soc.dbg_adr = 32'h24168; force soc.dbg_do = 32'h00021708; #1000;
force soc.dbg_adr = 32'h2416c; force soc.dbg_do = 32'h000216a4; #1000;
force soc.dbg_adr = 32'h24170; force soc.dbg_do = 32'h000216fc; #1000;
force soc.dbg_adr = 32'h24174; force soc.dbg_do = 32'h000216a4; #1000;
force soc.dbg_adr = 32'h24178; force soc.dbg_do = 32'h000216a4; #1000;
force soc.dbg_adr = 32'h2417c; force soc.dbg_do = 32'h000216f0; #1000;
force soc.dbg_adr = 32'h24180; force soc.dbg_do = 32'h000219dc; #1000;
force soc.dbg_adr = 32'h24184; force soc.dbg_do = 32'h00021738; #1000;
force soc.dbg_adr = 32'h24188; force soc.dbg_do = 32'h000219cc; #1000;
force soc.dbg_adr = 32'h2418c; force soc.dbg_do = 32'h00021738; #1000;
force soc.dbg_adr = 32'h24190; force soc.dbg_do = 32'h000219b0; #1000;
force soc.dbg_adr = 32'h24194; force soc.dbg_do = 32'h00021738; #1000;
force soc.dbg_adr = 32'h24198; force soc.dbg_do = 32'h00021738; #1000;
force soc.dbg_adr = 32'h2419c; force soc.dbg_do = 32'h00021738; #1000;
force soc.dbg_adr = 32'h241a0; force soc.dbg_do = 32'h00021738; #1000;
force soc.dbg_adr = 32'h241a4; force soc.dbg_do = 32'h00021738; #1000;
force soc.dbg_adr = 32'h241a8; force soc.dbg_do = 32'h00021738; #1000;
force soc.dbg_adr = 32'h241ac; force soc.dbg_do = 32'h00021738; #1000;
force soc.dbg_adr = 32'h241b0; force soc.dbg_do = 32'h0002172c; #1000;
force soc.dbg_adr = 32'h241b4; force soc.dbg_do = 32'h00021738; #1000;
force soc.dbg_adr = 32'h241b8; force soc.dbg_do = 32'h00021738; #1000;
force soc.dbg_adr = 32'h241bc; force soc.dbg_do = 32'h00021738; #1000;
force soc.dbg_adr = 32'h241c0; force soc.dbg_do = 32'h00021738; #1000;
force soc.dbg_adr = 32'h241c4; force soc.dbg_do = 32'h00021738; #1000;
force soc.dbg_adr = 32'h241c8; force soc.dbg_do = 32'h0002172c; #1000;
force soc.dbg_adr = 32'h241cc; force soc.dbg_do = 32'h00023900; #1000;
force soc.dbg_adr = 32'h241d0; force soc.dbg_do = 32'h0002381c; #1000;
force soc.dbg_adr = 32'h241d4; force soc.dbg_do = 32'h000237fc; #1000;
force soc.dbg_adr = 32'h241d8; force soc.dbg_do = 32'h0002381c; #1000;
force soc.dbg_adr = 32'h241dc; force soc.dbg_do = 32'h000238ec; #1000;
force soc.dbg_adr = 32'h241e0; force soc.dbg_do = 32'h0002381c; #1000;
force soc.dbg_adr = 32'h241e4; force soc.dbg_do = 32'h000237fc; #1000;
force soc.dbg_adr = 32'h241e8; force soc.dbg_do = 32'h00023900; #1000;
force soc.dbg_adr = 32'h241ec; force soc.dbg_do = 32'h00023900; #1000;
force soc.dbg_adr = 32'h241f0; force soc.dbg_do = 32'h000238ec; #1000;
force soc.dbg_adr = 32'h241f4; force soc.dbg_do = 32'h000237fc; #1000;
force soc.dbg_adr = 32'h241f8; force soc.dbg_do = 32'h00023828; #1000;
force soc.dbg_adr = 32'h241fc; force soc.dbg_do = 32'h00023828; #1000;
force soc.dbg_adr = 32'h24200; force soc.dbg_do = 32'h00023828; #1000;
force soc.dbg_adr = 32'h24204; force soc.dbg_do = 32'h000238ec; #1000;
force soc.dbg_adr = 32'h24208; force soc.dbg_do = 32'h02020100; #1000;
force soc.dbg_adr = 32'h2420c; force soc.dbg_do = 32'h03030303; #1000;
force soc.dbg_adr = 32'h24210; force soc.dbg_do = 32'h04040404; #1000;
force soc.dbg_adr = 32'h24214; force soc.dbg_do = 32'h04040404; #1000;
force soc.dbg_adr = 32'h24218; force soc.dbg_do = 32'h05050505; #1000;
force soc.dbg_adr = 32'h2421c; force soc.dbg_do = 32'h05050505; #1000;
force soc.dbg_adr = 32'h24220; force soc.dbg_do = 32'h05050505; #1000;
force soc.dbg_adr = 32'h24224; force soc.dbg_do = 32'h05050505; #1000;
force soc.dbg_adr = 32'h24228; force soc.dbg_do = 32'h06060606; #1000;
force soc.dbg_adr = 32'h2422c; force soc.dbg_do = 32'h06060606; #1000;
force soc.dbg_adr = 32'h24230; force soc.dbg_do = 32'h06060606; #1000;
force soc.dbg_adr = 32'h24234; force soc.dbg_do = 32'h06060606; #1000;
force soc.dbg_adr = 32'h24238; force soc.dbg_do = 32'h06060606; #1000;
force soc.dbg_adr = 32'h2423c; force soc.dbg_do = 32'h06060606; #1000;
force soc.dbg_adr = 32'h24240; force soc.dbg_do = 32'h06060606; #1000;
force soc.dbg_adr = 32'h24244; force soc.dbg_do = 32'h06060606; #1000;
force soc.dbg_adr = 32'h24248; force soc.dbg_do = 32'h07070707; #1000;
force soc.dbg_adr = 32'h2424c; force soc.dbg_do = 32'h07070707; #1000;
force soc.dbg_adr = 32'h24250; force soc.dbg_do = 32'h07070707; #1000;
force soc.dbg_adr = 32'h24254; force soc.dbg_do = 32'h07070707; #1000;
force soc.dbg_adr = 32'h24258; force soc.dbg_do = 32'h07070707; #1000;
force soc.dbg_adr = 32'h2425c; force soc.dbg_do = 32'h07070707; #1000;
force soc.dbg_adr = 32'h24260; force soc.dbg_do = 32'h07070707; #1000;
force soc.dbg_adr = 32'h24264; force soc.dbg_do = 32'h07070707; #1000;
force soc.dbg_adr = 32'h24268; force soc.dbg_do = 32'h07070707; #1000;
force soc.dbg_adr = 32'h2426c; force soc.dbg_do = 32'h07070707; #1000;
force soc.dbg_adr = 32'h24270; force soc.dbg_do = 32'h07070707; #1000;
force soc.dbg_adr = 32'h24274; force soc.dbg_do = 32'h07070707; #1000;
force soc.dbg_adr = 32'h24278; force soc.dbg_do = 32'h07070707; #1000;
force soc.dbg_adr = 32'h2427c; force soc.dbg_do = 32'h07070707; #1000;
force soc.dbg_adr = 32'h24280; force soc.dbg_do = 32'h07070707; #1000;
force soc.dbg_adr = 32'h24284; force soc.dbg_do = 32'h07070707; #1000;
force soc.dbg_adr = 32'h24288; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h2428c; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h24290; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h24294; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h24298; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h2429c; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242a0; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242a4; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242a8; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242ac; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242b0; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242b4; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242b8; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242bc; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242c0; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242c4; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242c8; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242cc; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242d0; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242d4; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242d8; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242dc; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242e0; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242e4; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242e8; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242ec; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242f0; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242f4; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242f8; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h242fc; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h24300; force soc.dbg_do = 32'h08080808; #1000;
force soc.dbg_adr = 32'h24304; force soc.dbg_do = 32'h08080808; #1000;

	release soc.cpu_n_reset;
	release soc.dbg_mem_op;
	release soc.dbg_wren;
	release soc.dbg_adr;
	release soc.dbg_do;
end

chaz #(
	.F_CLK(SIM_FCLK),
	.BAUD(SIM_BAUD)
) soc (
	.RESET(n_reset),
	.PICO_UART0_RX(rx),
	.PICO_UART0_TX(tx)
);

initial
begin
	$dumpfile(`VCD_OUTPUT);
	$dumpvars(3, t20_custom);
	#(40000000)
	$finish;
end

endmodule
