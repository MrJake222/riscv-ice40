../hazard3_config.vh