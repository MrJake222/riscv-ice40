../hazard3_width_const.vh