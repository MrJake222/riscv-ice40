parameter W_ADDR              = 32;
parameter W_DATA              = 32;
parameter NUM_IRQS            = 1;

module hazard3_noMAC (
	input wire                 clk,
	input wire                 clk_always_on,
	input wire                 rst_n,
	output wire                pwrup_req,
	input  wire                pwrup_ack,
	output wire                clk_en,
	output reg                 unblock_out,
	input  wire                unblock_in,
	output wire                bus_aph_req_i,
	output wire                bus_aph_panic_i, // e.g. branch mispredict + flush
	input  wire                bus_aph_ready_i,
	input  wire                bus_dph_ready_i,
	input  wire                bus_dph_err_i,
	output wire [W_ADDR-1:0]   bus_haddr_i,
	output wire [2:0]          bus_hsize_i,
	output wire                bus_priv_i,
	input  wire [W_DATA-1:0]   bus_rdata_i,
	output reg                 bus_aph_req_d,
	output wire                bus_aph_excl_d,
	input  wire                bus_aph_ready_d,
	input  wire                bus_dph_ready_d,
	input  wire                bus_dph_err_d,
	input  wire                bus_dph_exokay_d,
	output reg  [W_ADDR-1:0]   bus_haddr_d,
	output reg  [2:0]          bus_hsize_d,
	output reg                 bus_priv_d,
	output reg                 bus_hwrite_d,
	output reg  [W_DATA-1:0]   bus_wdata_d,
	input  wire [W_DATA-1:0]   bus_rdata_d,
	input  wire                dbg_req_halt,
	input  wire                dbg_req_halt_on_reset,
	input  wire                dbg_req_resume,
	output wire                dbg_halted,
	output wire                dbg_running,
	input  wire [W_DATA-1:0]   dbg_data0_rdata,
	output wire [W_DATA-1:0]   dbg_data0_wdata,
	output wire                dbg_data0_wen,
	input  wire [W_DATA-1:0]   dbg_instr_data,
	input  wire                dbg_instr_data_vld,
	output wire                dbg_instr_data_rdy,
	output wire                dbg_instr_caught_exception,
	output wire                dbg_instr_caught_ebreak,
	input  wire [NUM_IRQS-1:0] irq,       // -> mip.meip
	input  wire                soft_irq,  // -> mip.msip
	input  wire                timer_irq  // -> mip.mtip
);

hazard3_core #(
	.EXTENSION_M(0),
	.EXTENSION_A(0),
	.EXTENSION_C(0),
	.CSR_M_MANDATORY(0),
	.CSR_M_TRAP(0),
	.CSR_COUNTER(1)
) uut (
	.clk(clk),
	.clk_always_on(clk_always_on),
	.rst_n(rst_n),
	.pwrup_req(pwrup_req),
	.pwrup_ack(pwrup_ack),
	.clk_en(clk_en),
	.unblock_out(unblock_out),
	.unblock_in(unblock_in),
	.bus_aph_req_i(bus_aph_req_i),
	.bus_aph_panic_i(bus_aph_panic_i),
	.bus_aph_ready_i(bus_aph_ready_i),
	.bus_dph_ready_i(bus_dph_ready_i),
	.bus_dph_err_i(bus_dph_err_i),
	.bus_haddr_i(bus_haddr_i),
	.bus_hsize_i(bus_hsize_i),
	.bus_priv_i(bus_priv_i),
	.bus_rdata_i(bus_rdata_i),
	.bus_aph_req_d(bus_aph_req_d),
	.bus_aph_excl_d(bus_aph_excl_d),
	.bus_aph_ready_d(bus_aph_ready_d),
	.bus_dph_ready_d(bus_dph_ready_d),
	.bus_dph_err_d(bus_dph_err_d),
	.bus_dph_exokay_d(bus_dph_exokay_d),
	.bus_haddr_d(bus_haddr_d),
	.bus_hsize_d(bus_hsize_d),
	.bus_priv_d(bus_priv_d),
	.bus_hwrite_d(bus_hwrite_d),
	.bus_wdata_d(bus_wdata_d),
	.bus_rdata_d(bus_rdata_d),
	.dbg_req_halt(dbg_req_halt),
	.dbg_req_halt_on_reset(dbg_req_halt_on_reset),
	.dbg_req_resume(dbg_req_resume),
	.dbg_halted(dbg_halted),
	.dbg_running(dbg_running),
	.dbg_data0_rdata(dbg_data0_rdata),
	.dbg_data0_wdata(dbg_data0_wdata),
	.dbg_data0_wen(dbg_data0_wen),
	.dbg_instr_data(dbg_instr_data),
	.dbg_instr_data_vld(dbg_instr_data_vld),
	.dbg_instr_data_rdy(dbg_instr_data_rdy),
	.dbg_instr_caught_exception(dbg_instr_caught_exception),
	.dbg_instr_caught_ebreak(dbg_instr_caught_ebreak),
	.irq(irq),
	.soft_irq(soft_irq),
	.timer_irq(timer_irq)
);

endmodule
