../hazard3/hdl/hazard3_ops.vh